module top(
  input i_ce,
  input i_clk,
  input i_d1,
  input i_d2,
  input i_rst,
  output [23:0] io
  );
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_CE;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_I;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  wire [0:0] LIOB33_X0Y21_IOB_X0Y22_O;
  wire [0:0] LIOB33_X0Y23_IOB_X0Y23_O;
  wire [0:0] LIOB33_X0Y23_IOB_X0Y24_O;
  wire [0:0] LIOB33_X0Y25_IOB_X0Y25_O;
  wire [0:0] LIOB33_X0Y25_IOB_X0Y26_O;
  wire [0:0] LIOB33_X0Y27_IOB_X0Y27_O;
  wire [0:0] LIOB33_X0Y27_IOB_X0Y28_O;
  wire [0:0] LIOB33_X0Y29_IOB_X0Y29_O;
  wire [0:0] LIOB33_X0Y29_IOB_X0Y30_O;
  wire [0:0] LIOB33_X0Y31_IOB_X0Y31_O;
  wire [0:0] LIOB33_X0Y31_IOB_X0Y32_O;
  wire [0:0] LIOB33_X0Y33_IOB_X0Y33_O;
  wire [0:0] LIOB33_X0Y33_IOB_X0Y34_O;
  wire [0:0] LIOB33_X0Y35_IOB_X0Y35_O;
  wire [0:0] LIOB33_X0Y35_IOB_X0Y36_O;
  wire [0:0] LIOB33_X0Y37_IOB_X0Y37_O;
  wire [0:0] LIOB33_X0Y37_IOB_X0Y38_O;
  wire [0:0] LIOB33_X0Y39_IOB_X0Y39_O;
  wire [0:0] LIOB33_X0Y39_IOB_X0Y40_O;
  wire [0:0] LIOB33_X0Y41_IOB_X0Y41_O;
  wire [0:0] LIOB33_X0Y41_IOB_X0Y42_O;
  wire [0:0] LIOB33_X0Y43_IOB_X0Y43_O;
  wire [0:0] LIOB33_X0Y45_IOB_X0Y45_O;
  wire [0:0] LIOB33_X0Y45_IOB_X0Y46_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_CLK;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_D2;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_OCE;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_SR;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_CLK;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_D2;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_OCE;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_SR;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_CLK;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D2;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OCE;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_SR;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_CLK;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_D2;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_OCE;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_SR;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_CLK;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_D2;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_OCE;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_SR;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_TQ;
  wire [0:0] LIOI3_X0Y21_OLOGIC_X0Y22_CLK;
  wire [0:0] LIOI3_X0Y21_OLOGIC_X0Y22_D1;
  wire [0:0] LIOI3_X0Y21_OLOGIC_X0Y22_D2;
  wire [0:0] LIOI3_X0Y21_OLOGIC_X0Y22_OCE;
  wire [0:0] LIOI3_X0Y21_OLOGIC_X0Y22_OQ;
  wire [0:0] LIOI3_X0Y21_OLOGIC_X0Y22_SR;
  wire [0:0] LIOI3_X0Y21_OLOGIC_X0Y22_T1;
  wire [0:0] LIOI3_X0Y21_OLOGIC_X0Y22_TQ;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y23_CLK;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y23_D1;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y23_D2;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y23_OCE;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y23_OQ;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y23_SR;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y23_T1;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y23_TQ;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y24_CLK;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y24_D1;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y24_D2;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y24_OCE;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y24_OQ;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y24_SR;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y24_T1;
  wire [0:0] LIOI3_X0Y23_OLOGIC_X0Y24_TQ;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y25_CLK;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y25_D1;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y25_D2;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y25_OCE;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y25_OQ;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y25_SR;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y25_T1;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y25_TQ;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y26_CLK;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y26_D1;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y26_D2;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y26_OCE;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y26_OQ;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y26_SR;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y26_T1;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y26_TQ;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y27_CLK;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y27_D1;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y27_D2;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y27_OCE;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y27_OQ;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y27_SR;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y27_T1;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y27_TQ;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_CLK;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_D1;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_D2;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_OCE;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_OQ;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_SR;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_T1;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_TQ;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y29_CLK;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y29_D1;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y29_D2;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y29_OCE;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y29_OQ;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y29_SR;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y29_T1;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y29_TQ;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y30_CLK;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y30_D1;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y30_D2;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y30_OCE;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y30_OQ;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y30_SR;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y30_T1;
  wire [0:0] LIOI3_X0Y29_OLOGIC_X0Y30_TQ;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y33_CLK;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y33_D1;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y33_D2;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y33_OCE;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y33_OQ;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y33_SR;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y33_T1;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y33_TQ;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y34_CLK;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y34_D1;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y34_D2;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y34_OCE;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y34_OQ;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y34_SR;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y34_T1;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y34_TQ;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y35_CLK;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y35_D1;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y35_D2;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y35_OCE;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y35_OQ;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y35_SR;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y35_T1;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y35_TQ;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y36_CLK;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y36_D1;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y36_D2;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y36_OCE;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y36_OQ;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y36_SR;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y36_T1;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y36_TQ;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y39_CLK;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y39_D1;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y39_D2;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y39_OCE;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y39_OQ;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y39_SR;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y39_T1;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y39_TQ;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y40_CLK;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y40_D1;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y40_D2;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y40_OCE;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y40_OQ;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y40_SR;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y40_T1;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y40_TQ;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y41_CLK;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y41_D1;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y41_D2;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y41_OCE;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y41_OQ;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y41_SR;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y41_T1;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y41_TQ;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y42_CLK;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y42_D1;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y42_D2;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y42_OCE;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y42_OQ;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y42_SR;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y42_T1;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y42_TQ;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y45_CLK;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y45_D1;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y45_D2;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y45_OCE;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y45_OQ;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y45_SR;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y45_T1;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y45_TQ;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y46_CLK;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y46_D1;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y46_D2;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y46_OCE;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y46_OQ;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y46_SR;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y46_T1;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y46_TQ;
  wire [0:0] RIOB33_X43Y25_IOB_X1Y26_I;
  wire [0:0] RIOB33_X43Y43_IOB_X1Y43_I;
  wire [0:0] RIOB33_X43Y43_IOB_X1Y44_I;
  wire [0:0] RIOB33_X43Y45_IOB_X1Y45_I;
  wire [0:0] RIOB33_X43Y45_IOB_X1Y46_I;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_D;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_O;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_D;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_O;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_D;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_O;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y45_D;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y45_O;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y46_D;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y46_O;


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X43Y25_IOB_X1Y26_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y21_IOB_X0Y22_OBUF (
.I(LIOI3_X0Y21_OLOGIC_X0Y22_OQ),
.O(io[23])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y23_IOB_X0Y23_OBUF (
.I(LIOI3_X0Y23_OLOGIC_X0Y23_OQ),
.O(io[22])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y23_IOB_X0Y24_OBUF (
.I(LIOI3_X0Y23_OLOGIC_X0Y24_OQ),
.O(io[21])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y25_IOB_X0Y25_OBUF (
.I(LIOI3_X0Y25_OLOGIC_X0Y25_OQ),
.O(io[20])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y25_IOB_X0Y26_OBUF (
.I(LIOI3_X0Y25_OLOGIC_X0Y26_OQ),
.O(io[19])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y27_IOB_X0Y27_OBUF (
.I(LIOI3_X0Y27_OLOGIC_X0Y27_OQ),
.O(io[18])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y27_IOB_X0Y28_OBUF (
.I(LIOI3_X0Y27_OLOGIC_X0Y28_OQ),
.O(io[17])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y29_IOB_X0Y29_OBUF (
.I(LIOI3_X0Y29_OLOGIC_X0Y29_OQ),
.O(io[16])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y29_IOB_X0Y30_OBUF (
.I(LIOI3_X0Y29_OLOGIC_X0Y30_OQ),
.O(io[15])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y31_IOB_X0Y31_OBUF (
.I(LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_OQ),
.O(io[14])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y31_IOB_X0Y32_OBUF (
.I(LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_OQ),
.O(io[13])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y33_IOB_X0Y33_OBUF (
.I(LIOI3_X0Y33_OLOGIC_X0Y33_OQ),
.O(io[12])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y33_IOB_X0Y34_OBUF (
.I(LIOI3_X0Y33_OLOGIC_X0Y34_OQ),
.O(io[11])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y35_IOB_X0Y35_OBUF (
.I(LIOI3_X0Y35_OLOGIC_X0Y35_OQ),
.O(io[10])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y35_IOB_X0Y36_OBUF (
.I(LIOI3_X0Y35_OLOGIC_X0Y36_OQ),
.O(io[9])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y37_IOB_X0Y37_OBUF (
.I(LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_OQ),
.O(io[8])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y37_IOB_X0Y38_OBUF (
.I(LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_OQ),
.O(io[7])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y39_IOB_X0Y39_OBUF (
.I(LIOI3_X0Y39_OLOGIC_X0Y39_OQ),
.O(io[6])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y39_IOB_X0Y40_OBUF (
.I(LIOI3_X0Y39_OLOGIC_X0Y40_OQ),
.O(io[5])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y41_IOB_X0Y41_OBUF (
.I(LIOI3_X0Y41_OLOGIC_X0Y41_OQ),
.O(io[4])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y41_IOB_X0Y42_OBUF (
.I(LIOI3_X0Y41_OLOGIC_X0Y42_OQ),
.O(io[3])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y43_IOB_X0Y43_OBUF (
.I(LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ),
.O(io[2])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y45_IOB_X0Y45_OBUF (
.I(LIOI3_X0Y45_OLOGIC_X0Y45_OQ),
.O(io[1])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y45_IOB_X0Y46_OBUF (
.I(LIOI3_X0Y45_OLOGIC_X0Y46_OQ),
.O(io[0])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y21_OLOGIC_X0Y22_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y21_OLOGIC_X0Y22_OQ),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y23_OLOGIC_X0Y24_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y23_OLOGIC_X0Y24_OQ),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y23_OLOGIC_X0Y23_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y23_OLOGIC_X0Y23_OQ),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y25_OLOGIC_X0Y26_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y25_OLOGIC_X0Y26_OQ),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y25_OLOGIC_X0Y25_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y25_OLOGIC_X0Y25_OQ),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y27_OLOGIC_X0Y28_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y27_OLOGIC_X0Y28_OQ),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y27_OLOGIC_X0Y27_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y27_OLOGIC_X0Y27_OQ),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y29_OLOGIC_X0Y30_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y29_OLOGIC_X0Y30_OQ),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y29_OLOGIC_X0Y29_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y29_OLOGIC_X0Y29_OQ),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y33_OLOGIC_X0Y34_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y33_OLOGIC_X0Y34_OQ),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y33_OLOGIC_X0Y33_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y33_OLOGIC_X0Y33_OQ),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y35_OLOGIC_X0Y36_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y35_OLOGIC_X0Y36_OQ),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y35_OLOGIC_X0Y35_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y35_OLOGIC_X0Y35_OQ),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y39_OLOGIC_X0Y40_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y39_OLOGIC_X0Y40_OQ),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y39_OLOGIC_X0Y39_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y39_OLOGIC_X0Y39_OQ),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y41_OLOGIC_X0Y42_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y41_OLOGIC_X0Y42_OQ),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y41_OLOGIC_X0Y41_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y41_OLOGIC_X0Y41_OQ),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y45_OLOGIC_X0Y46_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y45_OLOGIC_X0Y46_OQ),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y45_OLOGIC_X0Y45_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_X0Y45_OLOGIC_X0Y45_OQ),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_OQ),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_OQ),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_OQ),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTFF" *)
  ODDR #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D1_INVERTED(1'b0),
    .IS_D2_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_ODDR_OQ (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D1(RIOB33_X43Y43_IOB_X1Y44_I),
.D2(RIOB33_X43Y43_IOB_X1Y43_I),
.Q(LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_OQ),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y25_IOB_X1Y26_IBUF (
.I(i_clk),
.O(RIOB33_X43Y25_IOB_X1Y26_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y43_IOB_X1Y43_IBUF (
.I(i_d2),
.O(RIOB33_X43Y43_IOB_X1Y43_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y43_IOB_X1Y44_IBUF (
.I(i_d1),
.O(RIOB33_X43Y43_IOB_X1Y44_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y45_IOB_X1Y45_IBUF (
.I(i_ce),
.O(RIOB33_X43Y45_IOB_X1Y45_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y45_IOB_X1Y46_IBUF (
.I(i_rst),
.O(RIOB33_X43Y45_IOB_X1Y46_I)
  );
  assign LIOI3_X0Y21_OLOGIC_X0Y22_TQ = LIOI3_X0Y21_OLOGIC_X0Y22_T1;
  assign LIOI3_X0Y23_OLOGIC_X0Y24_TQ = LIOI3_X0Y23_OLOGIC_X0Y24_T1;
  assign LIOI3_X0Y23_OLOGIC_X0Y23_TQ = LIOI3_X0Y23_OLOGIC_X0Y23_T1;
  assign LIOI3_X0Y25_OLOGIC_X0Y26_TQ = LIOI3_X0Y25_OLOGIC_X0Y26_T1;
  assign LIOI3_X0Y25_OLOGIC_X0Y25_TQ = LIOI3_X0Y25_OLOGIC_X0Y25_T1;
  assign LIOI3_X0Y27_OLOGIC_X0Y28_TQ = LIOI3_X0Y27_OLOGIC_X0Y28_T1;
  assign LIOI3_X0Y27_OLOGIC_X0Y27_TQ = LIOI3_X0Y27_OLOGIC_X0Y27_T1;
  assign LIOI3_X0Y29_OLOGIC_X0Y30_TQ = LIOI3_X0Y29_OLOGIC_X0Y30_T1;
  assign LIOI3_X0Y29_OLOGIC_X0Y29_TQ = LIOI3_X0Y29_OLOGIC_X0Y29_T1;
  assign LIOI3_X0Y33_OLOGIC_X0Y34_TQ = LIOI3_X0Y33_OLOGIC_X0Y34_T1;
  assign LIOI3_X0Y33_OLOGIC_X0Y33_TQ = LIOI3_X0Y33_OLOGIC_X0Y33_T1;
  assign LIOI3_X0Y35_OLOGIC_X0Y36_TQ = LIOI3_X0Y35_OLOGIC_X0Y36_T1;
  assign LIOI3_X0Y35_OLOGIC_X0Y35_TQ = LIOI3_X0Y35_OLOGIC_X0Y35_T1;
  assign LIOI3_X0Y39_OLOGIC_X0Y40_TQ = LIOI3_X0Y39_OLOGIC_X0Y40_T1;
  assign LIOI3_X0Y39_OLOGIC_X0Y39_TQ = LIOI3_X0Y39_OLOGIC_X0Y39_T1;
  assign LIOI3_X0Y41_OLOGIC_X0Y42_TQ = LIOI3_X0Y41_OLOGIC_X0Y42_T1;
  assign LIOI3_X0Y41_OLOGIC_X0Y41_TQ = LIOI3_X0Y41_OLOGIC_X0Y41_T1;
  assign LIOI3_X0Y45_OLOGIC_X0Y46_TQ = LIOI3_X0Y45_OLOGIC_X0Y46_T1;
  assign LIOI3_X0Y45_OLOGIC_X0Y45_TQ = LIOI3_X0Y45_OLOGIC_X0Y45_T1;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_TQ = LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_T1;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_TQ = LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_T1;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ = LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_TQ = LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_T1;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_TQ = LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_T1;
  assign RIOI3_X43Y25_ILOGIC_X1Y26_O = RIOI3_X43Y25_ILOGIC_X1Y26_D;
  assign RIOI3_X43Y45_ILOGIC_X1Y46_O = RIOI3_X43Y45_ILOGIC_X1Y46_D;
  assign RIOI3_X43Y45_ILOGIC_X1Y45_O = RIOI3_X43Y45_ILOGIC_X1Y45_D;
  assign RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_O = RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_D;
  assign RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_O = RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_D;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOB33_X0Y37_IOB_X0Y38_O = LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_OQ;
  assign LIOB33_X0Y37_IOB_X0Y37_O = LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_OQ;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_SR = 1'b0;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_SR = 1'b0;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_X0Y41_OLOGIC_X0Y42_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y41_OLOGIC_X0Y42_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y41_OLOGIC_X0Y42_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y41_OLOGIC_X0Y42_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y41_OLOGIC_X0Y42_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y41_OLOGIC_X0Y41_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOB33_X0Y41_IOB_X0Y42_O = LIOI3_X0Y41_OLOGIC_X0Y42_OQ;
  assign LIOB33_X0Y41_IOB_X0Y41_O = LIOI3_X0Y41_OLOGIC_X0Y41_OQ;
  assign LIOI3_X0Y41_OLOGIC_X0Y41_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y41_OLOGIC_X0Y41_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOB33_X0Y23_IOB_X0Y24_O = LIOI3_X0Y23_OLOGIC_X0Y24_OQ;
  assign LIOB33_X0Y23_IOB_X0Y23_O = LIOI3_X0Y23_OLOGIC_X0Y23_OQ;
  assign LIOI3_X0Y41_OLOGIC_X0Y41_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y41_OLOGIC_X0Y41_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y35_OLOGIC_X0Y36_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y35_OLOGIC_X0Y36_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y35_OLOGIC_X0Y36_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_X0Y35_OLOGIC_X0Y36_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y35_OLOGIC_X0Y36_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y35_OLOGIC_X0Y35_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y35_OLOGIC_X0Y35_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y35_OLOGIC_X0Y35_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOB33_X0Y45_IOB_X0Y46_O = LIOI3_X0Y45_OLOGIC_X0Y46_OQ;
  assign LIOB33_X0Y45_IOB_X0Y45_O = LIOI3_X0Y45_OLOGIC_X0Y45_OQ;
  assign LIOI3_X0Y35_OLOGIC_X0Y35_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOB33_X0Y27_IOB_X0Y28_O = LIOI3_X0Y27_OLOGIC_X0Y28_OQ;
  assign LIOB33_X0Y27_IOB_X0Y27_O = LIOI3_X0Y27_OLOGIC_X0Y27_OQ;
  assign LIOI3_X0Y35_OLOGIC_X0Y35_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y29_OLOGIC_X0Y30_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y29_OLOGIC_X0Y30_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
  assign LIOI3_X0Y29_OLOGIC_X0Y30_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_X0Y29_OLOGIC_X0Y30_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y29_OLOGIC_X0Y30_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y29_OLOGIC_X0Y29_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y29_OLOGIC_X0Y29_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y29_OLOGIC_X0Y29_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_X0Y29_OLOGIC_X0Y29_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y29_OLOGIC_X0Y29_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOB33_X0Y31_IOB_X0Y32_O = LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_OQ;
  assign LIOB33_X0Y31_IOB_X0Y31_O = LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y31_OQ;
  assign LIOI3_X0Y25_OLOGIC_X0Y26_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y25_OLOGIC_X0Y26_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y25_OLOGIC_X0Y26_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_X0Y25_OLOGIC_X0Y26_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y25_OLOGIC_X0Y26_SR = 1'b0;
  assign LIOI3_X0Y25_OLOGIC_X0Y25_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y25_OLOGIC_X0Y25_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y25_OLOGIC_X0Y25_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_X0Y25_OLOGIC_X0Y25_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y25_OLOGIC_X0Y25_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y21_OLOGIC_X0Y22_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y21_OLOGIC_X0Y22_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y21_OLOGIC_X0Y22_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOB33_X0Y35_IOB_X0Y36_O = LIOI3_X0Y35_OLOGIC_X0Y36_OQ;
  assign LIOB33_X0Y35_IOB_X0Y35_O = LIOI3_X0Y35_OLOGIC_X0Y35_OQ;
  assign LIOI3_X0Y21_OLOGIC_X0Y22_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y21_OLOGIC_X0Y22_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y45_OLOGIC_X0Y46_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y45_OLOGIC_X0Y46_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y45_OLOGIC_X0Y46_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_CE = 1'b1;
  assign LIOI3_X0Y45_OLOGIC_X0Y46_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y45_OLOGIC_X0Y46_SR = 1'b0;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOB33_X0Y39_IOB_X0Y40_O = LIOI3_X0Y39_OLOGIC_X0Y40_OQ;
  assign LIOB33_X0Y39_IOB_X0Y39_O = LIOI3_X0Y39_OLOGIC_X0Y39_OQ;
  assign LIOI3_X0Y45_OLOGIC_X0Y45_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign LIOB33_X0Y21_IOB_X0Y22_O = LIOI3_X0Y21_OLOGIC_X0Y22_OQ;
  assign LIOI3_X0Y45_OLOGIC_X0Y45_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y45_OLOGIC_X0Y45_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_X0Y45_OLOGIC_X0Y45_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y45_OLOGIC_X0Y45_SR = 1'b0;
  assign LIOI3_X0Y39_OLOGIC_X0Y40_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y39_OLOGIC_X0Y40_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y39_OLOGIC_X0Y40_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_X0Y39_OLOGIC_X0Y40_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y39_OLOGIC_X0Y40_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y39_OLOGIC_X0Y39_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y39_OLOGIC_X0Y39_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y39_OLOGIC_X0Y39_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOB33_X0Y43_IOB_X0Y43_O = LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ;
  assign LIOB33_X0Y25_IOB_X0Y26_O = LIOI3_X0Y25_OLOGIC_X0Y26_OQ;
  assign LIOB33_X0Y25_IOB_X0Y25_O = LIOI3_X0Y25_OLOGIC_X0Y25_OQ;
  assign LIOI3_X0Y39_OLOGIC_X0Y39_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y39_OLOGIC_X0Y39_SR = 1'b0;
  assign LIOI3_X0Y33_OLOGIC_X0Y34_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y33_OLOGIC_X0Y34_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y33_OLOGIC_X0Y34_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_X0Y33_OLOGIC_X0Y34_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y33_OLOGIC_X0Y34_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y33_OLOGIC_X0Y33_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y33_OLOGIC_X0Y33_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y33_OLOGIC_X0Y33_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_X0Y33_OLOGIC_X0Y33_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y33_OLOGIC_X0Y33_SR = 1'b0;
  assign LIOB33_X0Y29_IOB_X0Y30_O = LIOI3_X0Y29_OLOGIC_X0Y30_OQ;
  assign LIOB33_X0Y29_IOB_X0Y29_O = LIOI3_X0Y29_OLOGIC_X0Y29_OQ;
  assign LIOI3_X0Y27_OLOGIC_X0Y28_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y27_OLOGIC_X0Y28_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y27_OLOGIC_X0Y28_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_X0Y27_OLOGIC_X0Y28_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y27_OLOGIC_X0Y28_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y27_OLOGIC_X0Y27_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0 = RIOB33_X43Y25_IOB_X1Y26_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign LIOI3_X0Y27_OLOGIC_X0Y27_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y27_OLOGIC_X0Y27_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_X0Y27_OLOGIC_X0Y27_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y27_OLOGIC_X0Y27_SR = 1'b0;
  assign LIOI3_X0Y23_OLOGIC_X0Y24_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOB33_X0Y33_IOB_X0Y34_O = LIOI3_X0Y33_OLOGIC_X0Y34_OQ;
  assign LIOB33_X0Y33_IOB_X0Y33_O = LIOI3_X0Y33_OLOGIC_X0Y33_OQ;
  assign LIOI3_X0Y23_OLOGIC_X0Y24_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y23_OLOGIC_X0Y24_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_X0Y23_OLOGIC_X0Y24_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y23_OLOGIC_X0Y24_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y23_OLOGIC_X0Y23_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y23_OLOGIC_X0Y23_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOI3_X0Y23_OLOGIC_X0Y23_D2 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign LIOI3_X0Y23_OLOGIC_X0Y23_OCE = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y23_OLOGIC_X0Y23_SR = RIOB33_X43Y45_IOB_X1Y46_I;
endmodule
