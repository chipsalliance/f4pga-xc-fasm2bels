module top(
  input clk,
  output [3:0] led,
  output tx
  );
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR0;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR1;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR10;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR11;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR12;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR13;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR2;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR3;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR4;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR5;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR6;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR7;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR8;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR9;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRATIEHIGH0;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRATIEHIGH1;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBTIEHIGH0;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBTIEHIGH1;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR0;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR1;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR10;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR11;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR12;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR13;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR2;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR3;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR4;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR5;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR6;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR7;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR8;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR9;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI0;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI1;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI10;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI11;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI12;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI13;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI14;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI15;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI2;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI3;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI4;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI5;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI6;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI7;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI8;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIADI9;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI0;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI1;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI10;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI11;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI12;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI13;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI14;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI15;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI2;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI3;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI4;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI5;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI6;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI7;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI8;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI9;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIPADIP0;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIPADIP1;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIPBDIP0;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DIPBDIP1;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO0;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO1;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO10;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO11;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO12;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO13;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO14;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO15;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO16;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO17;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO18;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO19;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO2;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO20;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO21;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO22;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO23;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO24;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO25;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO26;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO27;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO28;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO29;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO3;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO30;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO31;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO4;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO5;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO6;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO7;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO8;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DO9;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DOP0;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DOP1;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DOP2;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_DOP3;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_RDCLK;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_RDEN;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_RDRCLK;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_REGCE;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_REGCEB;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_REGCLKB;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_RST;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_RSTRAMB;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_RSTREG;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_RSTREGB;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_WEA0;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_WEA1;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_WEA2;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_WEA3;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE0;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE1;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE2;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE3;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE4;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE5;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE6;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE7;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_WRCLK;
  wire [0:0] BRAM_L_X44Y95_RAMB18_X2Y38_WREN;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_A;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_A1;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_A2;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_A3;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_A4;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_A5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_A5Q;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_A6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_AMUX;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_AO5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_AO6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_A_CY;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_A_XOR;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_B;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_B1;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_B2;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_B3;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_B4;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_B5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_B6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_BO5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_BO6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_B_CY;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_B_XOR;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_C;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_C1;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_C2;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_C3;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_C4;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_C5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_C6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_CE;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_CLK;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_CO5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_CO6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_C_CY;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_C_XOR;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_D;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_D1;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_D2;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_D3;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_D4;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_D5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_D6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_DO5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_DO6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_D_CY;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_D_XOR;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X68Y101_SR;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_A;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_A1;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_A2;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_A3;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_A4;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_A5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_A5Q;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_A6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_AMUX;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_AO5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_AO6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_AQ;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_AX;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_A_CY;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_A_XOR;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_B;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_B1;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_B2;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_B3;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_B4;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_B5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_B6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_BMUX;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_BO5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_BO6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_BQ;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_BX;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_B_CY;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_B_XOR;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_C;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_C1;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_C2;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_C3;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_C4;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_C5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_C5Q;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_C6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_CE;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_CLK;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_CMUX;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_CO5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_CO6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_CQ;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_CX;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_C_CY;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_C_XOR;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_D;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_D1;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_D2;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_D3;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_D4;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_D5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_D5Q;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_D6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_DMUX;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_DO5;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_DO6;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_DX;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_D_CY;
  wire [0:0] CLBLL_L_X42Y101_SLICE_X69Y101_D_XOR;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_A;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_A1;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_A2;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_A3;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_A4;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_A5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_A6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_AMUX;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_AO5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_AO6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_A_CY;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_A_XOR;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_B;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_B1;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_B2;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_B3;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_B4;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_B5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_B6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_BMUX;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_BO5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_BO6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_BQ;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_B_CY;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_B_XOR;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_C;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_C1;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_C2;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_C3;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_C4;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_C5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_C6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_CE;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_CLK;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_CMUX;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_CO5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_CO6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_C_CY;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_C_XOR;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_D;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_D1;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_D2;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_D3;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_D4;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_D5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_D6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_DMUX;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_DO5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_DO6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_D_CY;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_D_XOR;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X68Y102_SR;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_A;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_A1;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_A2;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_A3;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_A4;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_A5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_A5Q;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_A6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_AMUX;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_AO5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_AO6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_AQ;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_AX;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_A_CY;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_A_XOR;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_B;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_B1;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_B2;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_B3;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_B4;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_B5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_B6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_BMUX;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_BO5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_BO6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_B_CY;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_B_XOR;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_C;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_C1;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_C2;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_C3;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_C4;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_C5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_C5Q;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_C6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_CE;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_CLK;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_CMUX;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_CO5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_CO6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_CQ;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_CX;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_C_CY;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_C_XOR;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_D;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_D1;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_D2;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_D3;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_D4;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_D5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_D5Q;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_D6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_DMUX;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_DO5;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_DO6;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_DQ;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_DX;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_D_CY;
  wire [0:0] CLBLL_L_X42Y102_SLICE_X69Y102_D_XOR;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_A;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_A1;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_A2;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_A3;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_A4;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_A5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_A6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_AMUX;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_AO5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_AO6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_A_CY;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_A_XOR;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_B;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_B1;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_B2;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_B3;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_B4;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_B5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_B6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_BMUX;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_BO6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_BQ;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_BX;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_B_CY;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_B_XOR;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_C;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_C1;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_C2;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_C3;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_C4;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_C5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_C6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_CE;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_CLK;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_CMUX;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_CO5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_CO6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_CQ;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_CX;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_C_CY;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_C_XOR;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_D;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_D1;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_D2;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_D3;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_D4;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_D5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_D6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_DMUX;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_DO5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_DO6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_DQ;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_DX;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_D_CY;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X68Y103_D_XOR;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_A;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_A1;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_A2;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_A3;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_A4;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_A5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_A6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_AMUX;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_AO5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_AO6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_AX;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_A_CY;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_A_XOR;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_B;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_B1;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_B2;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_B3;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_B4;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_B5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_B6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_BMUX;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_BO5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_BO6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_BQ;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_BX;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_B_CY;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_B_XOR;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_C;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_C1;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_C2;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_C3;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_C4;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_C5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_C6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_CE;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_CLK;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_CMUX;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_CO5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_CO6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_COUT;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_CX;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_C_CY;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_C_XOR;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_D;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_D1;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_D2;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_D3;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_D4;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_D5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_D6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_DMUX;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_DO5;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_DO6;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_DX;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_D_CY;
  wire [0:0] CLBLL_L_X42Y103_SLICE_X69Y103_D_XOR;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_A;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_A1;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_A2;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_A3;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_A4;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_A5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_A6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_AMUX;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_AO5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_AO6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_A_CY;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_A_XOR;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_B;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_B1;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_B2;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_B3;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_B4;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_B5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_B6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_BMUX;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_BO5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_BO6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_B_CY;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_B_XOR;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_C;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_C1;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_C2;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_C3;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_C4;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_C5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_C6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_CE;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_CLK;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_CMUX;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_CO5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_CO6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_C_CY;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_C_XOR;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_D;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_D1;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_D2;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_D3;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_D4;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_D5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_D6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_DMUX;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_DO5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_DO6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_DX;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_D_CY;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X68Y104_D_XOR;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_A;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_A1;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_A2;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_A3;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_A4;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_A5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_A6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_AMUX;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_AO5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_AO6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_AQ;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_AX;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_A_CY;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_A_XOR;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_B;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_B1;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_B2;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_B3;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_B4;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_B5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_B6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_BMUX;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_BO5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_BO6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_BQ;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_BX;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_B_CY;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_B_XOR;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_C;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_C1;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_C2;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_C3;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_C4;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_C5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_C6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_CE;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_CIN;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_CLK;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_CMUX;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_CO5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_CO6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_COUT;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_CQ;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_CX;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_C_CY;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_C_XOR;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_D;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_D1;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_D2;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_D3;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_D4;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_D5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_D6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_DMUX;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_DO5;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_DO6;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_DX;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_D_XOR;
  wire [0:0] CLBLL_L_X42Y104_SLICE_X69Y104_SR;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_A;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_A1;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_A2;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_A3;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_A4;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_A5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_A6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_AMUX;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_AO5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_AO6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_A_CY;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_A_XOR;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_B;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_B1;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_B2;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_B3;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_B4;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_B5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_B6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_BMUX;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_BO5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_BO6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_B_CY;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_B_XOR;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_C;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_C1;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_C2;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_C3;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_C4;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_C5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_C6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_CE;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_CLK;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_CMUX;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_CO5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_CO6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_CQ;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_CX;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_C_CY;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_C_XOR;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_D;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_D1;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_D2;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_D3;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_D4;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_D5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_D6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_DMUX;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_DO5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_DO6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_D_CY;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X68Y105_D_XOR;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_A;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_A1;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_A2;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_A3;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_A4;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_A5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_A5Q;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_A6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_AMUX;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_AO5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_AO6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_AQ;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_AX;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_A_CY;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_A_XOR;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_B;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_B1;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_B2;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_B3;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_B4;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_B5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_B6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_BMUX;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_BO5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_BO6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_B_CY;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_B_XOR;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_C;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_C1;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_C2;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_C3;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_C4;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_C5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_C6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_CE;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_CLK;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_CMUX;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_CO5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_CO6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_C_CY;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_C_XOR;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_D;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_D1;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_D2;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_D3;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_D4;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_D5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_D6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_DMUX;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_DO5;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_DO6;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_D_CY;
  wire [0:0] CLBLL_L_X42Y105_SLICE_X69Y105_D_XOR;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_A;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_A1;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_A2;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_A3;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_A4;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_A5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_A5Q;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_A6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_AMUX;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_AO5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_AO6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_AQ;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_AX;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_A_CY;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_A_XOR;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_B;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_B1;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_B2;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_B3;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_B4;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_B5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_B6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_BMUX;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_BO5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_BO6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_B_CY;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_B_XOR;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_C;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_C1;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_C2;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_C3;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_C4;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_C5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_C6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_CE;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_CLK;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_CMUX;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_CO5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_CO6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_C_CY;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_C_XOR;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_D;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_D1;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_D2;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_D3;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_D4;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_D5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_D6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_DMUX;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_DO5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_DO6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_D_CY;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X68Y106_D_XOR;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_A;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_A1;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_A2;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_A3;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_A4;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_A5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_A6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_AMUX;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_AO5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_AO6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_A_CY;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_A_XOR;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_B;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_B1;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_B2;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_B3;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_B4;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_B5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_B6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_BMUX;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_BO5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_BO6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_B_CY;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_B_XOR;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_C;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_C1;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_C2;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_C3;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_C4;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_C5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_C6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_CE;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_CLK;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_CMUX;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_CO5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_CO6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_CQ;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_CX;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_C_CY;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_C_XOR;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_D;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_D1;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_D2;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_D3;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_D4;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_D5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_D6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_DMUX;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_DO5;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_DO6;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_D_CY;
  wire [0:0] CLBLL_L_X42Y106_SLICE_X69Y106_D_XOR;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_A;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_A1;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_A2;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_A3;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_A4;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_A5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_A6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_AMUX;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_AO5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_AO6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_A_CY;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_A_XOR;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_B;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_B1;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_B2;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_B3;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_B4;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_B5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_B6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_BMUX;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_BO5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_BO6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_BQ;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_BX;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_B_CY;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_B_XOR;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_C;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_C1;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_C2;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_C3;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_C4;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_C5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_C6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_CE;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_CLK;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_CMUX;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_CO5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_CO6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_C_CY;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_C_XOR;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_D;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_D1;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_D2;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_D3;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_D4;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_D5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_D6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_DMUX;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_DO5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_D_CY;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X68Y107_D_XOR;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_A;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_A1;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_A2;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_A3;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_A4;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_A5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_A5Q;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_A6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_AMUX;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_AO5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_AO6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_AQ;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_AX;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_A_CY;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_A_XOR;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_B;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_B1;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_B2;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_B3;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_B4;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_B5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_B5Q;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_B6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_BMUX;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_BO5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_BO6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_BQ;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_BX;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_B_CY;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_B_XOR;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_C;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_C1;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_C2;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_C3;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_C4;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_C5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_C5Q;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_C6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_CE;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_CLK;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_CMUX;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_CO5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_CO6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_CQ;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_CX;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_C_CY;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_C_XOR;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_D;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_D1;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_D2;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_D3;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_D4;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_D5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_D5Q;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_D6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_DMUX;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_DO5;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_DO6;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_DQ;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_DX;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_D_CY;
  wire [0:0] CLBLL_L_X42Y107_SLICE_X69Y107_D_XOR;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_A;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_A1;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_A2;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_A3;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_A4;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_A5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_A6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_AMUX;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_AO5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_AO6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_A_CY;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_A_XOR;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_B;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_B1;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_B2;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_B3;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_B4;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_B5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_B6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_BMUX;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_BO5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_BO6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_B_CY;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_B_XOR;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_C;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_C1;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_C2;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_C3;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_C4;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_C5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_C5Q;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_C6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_CE;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_CLK;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_CMUX;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_CO5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_CO6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_C_CY;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_C_XOR;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_D;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_D1;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_D2;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_D3;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_D4;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_D5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_D6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_DMUX;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_DO5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_DO6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_D_CY;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_D_XOR;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X68Y108_SR;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_A;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_A1;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_A2;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_A3;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_A4;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_A5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_A5Q;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_A6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_AMUX;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_AO5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_AO6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_AQ;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_AX;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_A_CY;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_A_XOR;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_B;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_B1;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_B2;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_B3;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_B4;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_B5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_B6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_BMUX;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_BO5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_BO6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_B_CY;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_B_XOR;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_C;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_C1;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_C2;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_C3;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_C4;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_C5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_C6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_CE;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_CLK;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_CMUX;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_CO5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_CO6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_C_CY;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_C_XOR;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_D;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_D1;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_D2;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_D3;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_D4;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_D5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_D5Q;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_D6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_DMUX;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_DO5;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_DO6;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_DQ;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_DX;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_D_CY;
  wire [0:0] CLBLL_L_X42Y108_SLICE_X69Y108_D_XOR;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_A;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_A1;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_A2;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_A3;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_A4;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_A5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_A6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_AMUX;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_AO5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_AO6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_A_CY;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_A_XOR;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_B;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_B1;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_B2;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_B3;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_B4;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_B5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_B6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_BMUX;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_BO5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_BO6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_B_CY;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_B_XOR;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_C;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_C1;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_C2;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_C3;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_C4;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_C5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_C6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_CLK;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_CMUX;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_CO5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_CO6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_C_CY;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_C_XOR;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_D;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_D1;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_D2;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_D3;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_D4;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_D5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_D5Q;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_D6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_DMUX;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_DO5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_DO6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_DQ;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_DX;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_D_CY;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_D_XOR;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X68Y109_SR;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_A;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_A1;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_A2;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_A3;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_A4;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_A5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_A6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_AMUX;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_AO5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_AO6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_A_CY;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_A_XOR;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_B;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_B1;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_B2;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_B3;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_B4;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_B5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_B6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_BMUX;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_BO5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_BO6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_B_CY;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_B_XOR;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_C;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_C1;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_C2;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_C3;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_C4;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_C5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_C6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_CE;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_CLK;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_CMUX;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_CO5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_CO6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_C_CY;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_C_XOR;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_D;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_D1;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_D2;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_D3;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_D4;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_D5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_D6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_DO5;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_DO6;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_DQ;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_D_CY;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_D_XOR;
  wire [0:0] CLBLL_L_X42Y109_SLICE_X69Y109_SR;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_A;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_A1;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_A2;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_A3;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_A4;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_A5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_A6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_AMUX;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_AO5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_AO6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_A_CY;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_A_XOR;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_B;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_B1;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_B2;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_B3;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_B4;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_B5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_B6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_BMUX;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_BO5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_BO6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_B_CY;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_B_XOR;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_C;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_C1;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_C2;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_C3;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_C4;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_C5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_C5Q;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_C6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_CE;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_CLK;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_CMUX;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_CO5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_CO6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_C_CY;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_C_XOR;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_D;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_D1;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_D2;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_D3;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_D4;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_D5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_D6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_DMUX;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_DO5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_DO6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_D_CY;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_D_XOR;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X68Y110_SR;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_A;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_A1;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_A2;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_A3;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_A4;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_A5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_A6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_AMUX;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_AO5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_AO6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_AQ;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_AX;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_A_CY;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_A_XOR;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_B;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_B1;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_B2;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_B3;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_B4;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_B5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_B6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_BMUX;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_BO5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_BO6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_BX;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_B_CY;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_B_XOR;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_C;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_C1;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_C2;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_C3;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_C4;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_C5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_C5Q;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_C6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_CLK;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_CMUX;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_CO5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_CO6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_C_CY;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_C_XOR;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_D;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_D1;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_D2;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_D3;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_D4;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_D5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_D6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_DMUX;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_DO5;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_DO6;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_D_CY;
  wire [0:0] CLBLL_L_X42Y110_SLICE_X69Y110_D_XOR;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_A;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_A1;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_A2;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_A3;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_A4;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_A5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_A5Q;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_A6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_AMUX;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_AO5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_AO6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_AQ;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_AX;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_A_CY;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_A_XOR;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_B;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_B1;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_B2;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_B3;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_B4;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_B5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_B5Q;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_B6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_BMUX;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_BO5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_BO6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_BQ;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_BX;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_B_CY;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_B_XOR;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_C;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_C1;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_C2;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_C3;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_C4;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_C5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_C5Q;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_C6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_CE;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_CLK;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_CMUX;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_CO5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_CO6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_CQ;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_CX;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_C_CY;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_C_XOR;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_D;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_D1;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_D2;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_D3;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_D4;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_D5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_D5Q;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_D6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_DMUX;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_DO5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_DO6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_DQ;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_DX;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_D_CY;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X68Y111_D_XOR;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_A;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_A1;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_A2;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_A3;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_A4;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_A5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_A5Q;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_A6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_AMUX;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_AO5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_AO6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_AQ;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_AX;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_A_CY;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_A_XOR;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_B;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_B1;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_B2;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_B3;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_B4;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_B5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_B6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_BO5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_BO6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_BQ;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_BX;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_B_CY;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_B_XOR;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_C;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_C1;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_C2;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_C3;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_C4;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_C5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_C6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_CE;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_CLK;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_CMUX;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_CO5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_CO6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_C_CY;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_C_XOR;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_D;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_D1;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_D2;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_D3;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_D4;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_D5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_D5Q;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_D6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_DMUX;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_DO5;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_DO6;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_DQ;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_DX;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_D_CY;
  wire [0:0] CLBLL_L_X42Y111_SLICE_X69Y111_D_XOR;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_A;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_A1;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_A2;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_A3;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_A4;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_A5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_A5Q;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_A6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_AMUX;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_AO5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_AO6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_AQ;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_AX;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_A_CY;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_A_XOR;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_B;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_B1;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_B2;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_B3;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_B4;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_B5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_B5Q;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_B6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_BMUX;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_BO5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_BO6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_BQ;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_BX;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_B_CY;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_B_XOR;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_C;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_C1;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_C2;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_C3;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_C4;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_C5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_C5Q;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_C6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_CE;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_CLK;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_CMUX;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_CO5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_CO6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_CQ;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_CX;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_C_CY;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_C_XOR;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_D;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_D1;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_D2;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_D3;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_D4;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_D5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_D5Q;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_D6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_DMUX;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_DO5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_DO6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_DQ;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_DX;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_D_CY;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X68Y112_D_XOR;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_A;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_A1;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_A2;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_A3;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_A4;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_A5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_A6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_AMUX;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_AO5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_AO6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_A_CY;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_A_XOR;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_B;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_B1;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_B2;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_B3;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_B4;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_B5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_B6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_BMUX;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_BO5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_BO6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_BQ;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_BX;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_B_CY;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_B_XOR;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_C;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_C1;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_C2;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_C3;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_C4;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_C5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_C5Q;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_C6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_CLK;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_CMUX;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_CO5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_CO6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_C_CY;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_C_XOR;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_D;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_D1;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_D2;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_D3;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_D4;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_D5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_D6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_DMUX;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_DO5;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_DO6;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_DQ;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_DX;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_D_CY;
  wire [0:0] CLBLL_L_X42Y112_SLICE_X69Y112_D_XOR;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_A;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_A1;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_A2;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_A3;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_A4;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_A5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_A6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_AO5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_AO6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_A_CY;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_A_XOR;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_B;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_B1;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_B2;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_B3;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_B4;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_B5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_B6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_BO5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_BO6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_B_CY;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_B_XOR;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_C;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_C1;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_C2;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_C3;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_C4;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_C5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_C6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_CE;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_CLK;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_CO5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_CO6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_C_CY;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_C_XOR;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_D;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_D1;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_D2;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_D3;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_D4;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_D5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_D5Q;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_D6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_DMUX;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_DO5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_DO6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_DX;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_D_CY;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_D_XOR;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X68Y113_SR;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_A;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_A1;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_A2;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_A3;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_A4;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_A5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_A5Q;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_A6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_AMUX;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_AO5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_AO6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_AQ;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_AX;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_A_CY;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_A_XOR;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_B;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_B1;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_B2;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_B3;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_B4;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_B5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_B5Q;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_B6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_BMUX;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_BO5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_BO6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_BQ;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_BX;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_B_CY;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_B_XOR;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_C;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_C1;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_C2;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_C3;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_C4;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_C5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_C5Q;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_C6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_CE;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_CLK;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_CMUX;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_CO5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_CO6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_CQ;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_CX;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_C_CY;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_C_XOR;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_D;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_D1;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_D2;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_D3;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_D4;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_D5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_D5Q;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_D6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_DMUX;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_DO5;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_DO6;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_DQ;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_DX;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_D_CY;
  wire [0:0] CLBLL_L_X42Y113_SLICE_X69Y113_D_XOR;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_A;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_A1;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_A2;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_A3;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_A4;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_A5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_A6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_AO5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_AO6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_A_CY;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_A_XOR;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_B;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_B1;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_B2;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_B3;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_B4;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_B5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_B6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_BO5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_BO6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_B_CY;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_B_XOR;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_C;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_C1;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_C2;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_C3;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_C4;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_C5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_C6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_CO5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_CO6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_C_CY;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_C_XOR;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_D;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_D1;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_D2;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_D3;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_D4;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_D5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_D6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_DO5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_DO6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_D_CY;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X68Y118_D_XOR;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_A;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_A1;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_A2;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_A3;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_A4;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_A5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_A5Q;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_A6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_AMUX;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_AO5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_AO6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_AQ;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_AX;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_A_CY;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_A_XOR;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_B;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_B1;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_B2;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_B3;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_B4;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_B5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_B5Q;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_B6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_BMUX;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_BO5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_BO6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_BQ;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_BX;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_B_CY;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_B_XOR;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_C;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_C1;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_C2;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_C3;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_C4;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_C5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_C5Q;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_C6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_CE;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_CLK;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_CMUX;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_CO5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_CO6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_CQ;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_CX;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_C_CY;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_C_XOR;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_D;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_D1;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_D2;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_D3;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_D4;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_D5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_D5Q;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_D6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_DMUX;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_DO5;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_DO6;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_DQ;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_DX;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_D_CY;
  wire [0:0] CLBLL_L_X42Y118_SLICE_X69Y118_D_XOR;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_A;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_A1;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_A2;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_A3;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_A4;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_A5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_A6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_AO5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_AO6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_AX;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_A_CY;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_A_XOR;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_B;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_B1;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_B2;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_B3;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_B4;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_B5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_B6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_BMUX;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_BO5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_BO6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_BX;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_B_CY;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_B_XOR;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_C;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_C1;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_C2;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_C3;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_C4;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_C5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_C6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_CMUX;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_CO5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_CO6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_COUT;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_CX;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_C_CY;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_C_XOR;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_D;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_D1;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_D2;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_D3;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_D4;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_D5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_D6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_DMUX;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_DO5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_DO6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_DX;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_D_CY;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X68Y43_D_XOR;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_A;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_A1;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_A2;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_A3;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_A4;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_A5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_A6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_AO5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_AO6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_A_CY;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_A_XOR;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_B;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_B1;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_B2;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_B3;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_B4;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_B5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_B6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_BO5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_BO6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_B_CY;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_B_XOR;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_C;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_C1;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_C2;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_C3;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_C4;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_C5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_C6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_CO5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_CO6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_C_CY;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_C_XOR;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_D;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_D1;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_D2;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_D3;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_D4;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_D5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_D6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_DO5;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_DO6;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_D_CY;
  wire [0:0] CLBLL_L_X42Y43_SLICE_X69Y43_D_XOR;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_A;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_A1;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_A2;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_A3;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_A4;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_A5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_A5Q;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_A6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_AMUX;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_AO5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_AO6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_AQ;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_AX;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_A_CY;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_A_XOR;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_B;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_B1;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_B2;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_B3;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_B4;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_B5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_B5Q;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_B6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_BMUX;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_BO5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_BO6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_BQ;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_BX;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_B_CY;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_B_XOR;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_C;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_C1;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_C2;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_C3;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_C4;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_C5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_C5Q;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_C6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_CE;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_CLK;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_CMUX;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_CO5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_CO6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_CQ;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_CX;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_C_CY;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_C_XOR;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_D;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_D1;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_D2;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_D3;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_D4;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_D5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_D5Q;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_D6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_DMUX;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_DO5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_DO6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_DQ;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_DX;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_D_CY;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X68Y68_D_XOR;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_A;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_A1;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_A2;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_A3;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_A4;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_A5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_A6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_AO5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_AO6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_A_CY;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_A_XOR;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_B;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_B1;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_B2;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_B3;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_B4;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_B5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_B6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_BO5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_BO6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_B_CY;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_B_XOR;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_C;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_C1;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_C2;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_C3;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_C4;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_C5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_C6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_CO5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_CO6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_C_CY;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_C_XOR;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_D;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_D1;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_D2;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_D3;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_D4;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_D5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_D6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_DO5;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_DO6;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_D_CY;
  wire [0:0] CLBLL_L_X42Y68_SLICE_X69Y68_D_XOR;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_A;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_A1;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_A2;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_A3;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_A4;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_A5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_A6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_AMUX;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_AO5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_AO6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_AQ;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_AX;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_A_CY;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_A_XOR;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_B;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_B1;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_B2;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_B3;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_B4;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_B5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_B6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_BMUX;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_BO5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_BO6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_BQ;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_BX;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_B_CY;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_B_XOR;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_C;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_C1;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_C2;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_C3;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_C4;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_C5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_C6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_CLK;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_CMUX;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_CO5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_CO6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_COUT;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_CQ;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_CX;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_C_CY;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_C_XOR;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_D;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_D1;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_D2;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_D3;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_D4;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_D5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_D6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_DMUX;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_DO5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_DO6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_DQ;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_DX;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_D_CY;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_D_XOR;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X68Y69_SR;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_A;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_A1;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_A2;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_A3;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_A4;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_A5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_A6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_AO5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_AO6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_A_CY;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_A_XOR;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_B;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_B1;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_B2;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_B3;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_B4;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_B5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_B6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_BO5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_BO6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_B_CY;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_B_XOR;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_C;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_C1;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_C2;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_C3;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_C4;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_C5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_C6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_CMUX;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_CO5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_CO6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_C_CY;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_C_XOR;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_D;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_D1;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_D2;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_D3;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_D4;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_D5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_D6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_DO5;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_DO6;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_D_CY;
  wire [0:0] CLBLL_L_X42Y69_SLICE_X69Y69_D_XOR;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_A;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_A1;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_A2;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_A3;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_A4;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_A5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_A6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_AMUX;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_AO5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_AO6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_AQ;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_AX;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_A_CY;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_A_XOR;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_B;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_B1;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_B2;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_B3;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_B4;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_B5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_B6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_BMUX;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_BO5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_BO6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_BQ;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_BX;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_B_CY;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_B_XOR;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_C;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_C1;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_C2;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_C3;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_C4;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_C5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_C6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_CIN;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_CLK;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_CMUX;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_CO5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_CO6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_COUT;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_CX;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_C_CY;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_C_XOR;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_D;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_D1;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_D2;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_D3;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_D4;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_D5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_D6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_DMUX;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_DO5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_DO6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_DQ;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_DX;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X68Y70_D_XOR;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_A;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_A1;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_A2;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_A3;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_A4;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_A5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_A6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_AO5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_AO6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_A_CY;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_A_XOR;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_B;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_B1;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_B2;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_B3;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_B4;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_B5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_B6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_BO5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_BO6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_B_CY;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_B_XOR;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_C;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_C1;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_C2;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_C3;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_C4;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_C5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_C6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_CO5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_CO6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_C_CY;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_C_XOR;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_D;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_D1;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_D2;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_D3;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_D4;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_D5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_D6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_DO5;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_DO6;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_D_CY;
  wire [0:0] CLBLL_L_X42Y70_SLICE_X69Y70_D_XOR;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_A;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_A1;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_A2;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_A3;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_A4;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_A5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_A6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_AMUX;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_AO5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_AO6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_A_CY;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_A_XOR;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_B;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_B1;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_B2;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_B3;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_B4;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_B5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_B5Q;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_B6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_BMUX;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_BO5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_BO6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_BQ;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_BX;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_B_CY;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_B_XOR;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_C;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_C1;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_C2;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_C3;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_C4;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_C5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_C6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_CLK;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_CMUX;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_CO5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_CO6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_C_CY;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_C_XOR;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_D;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_D1;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_D2;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_D3;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_D4;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_D5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_D6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_DMUX;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_DO5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_DO6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_D_CY;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_D_XOR;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X68Y71_SR;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_A;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_A1;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_A2;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_A3;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_A4;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_A5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_A6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_AO5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_AO6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_A_CY;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_A_XOR;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_B;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_B1;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_B2;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_B3;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_B4;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_B5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_B6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_BO5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_BO6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_B_CY;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_B_XOR;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_C;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_C1;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_C2;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_C3;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_C4;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_C5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_C6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_CO5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_CO6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_C_CY;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_C_XOR;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_D;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_D1;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_D2;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_D3;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_D4;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_D5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_D6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_DO5;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_DO6;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_D_CY;
  wire [0:0] CLBLL_L_X42Y71_SLICE_X69Y71_D_XOR;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_A;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_A1;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_A2;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_A3;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_A4;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_A5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_A6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_AO5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_AO6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_A_CY;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_A_XOR;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_B;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_B1;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_B2;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_B3;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_B4;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_B5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_B6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_BO5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_BO6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_B_CY;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_B_XOR;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_C;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_C1;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_C2;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_C3;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_C4;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_C5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_C6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_CO5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_CO6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_C_CY;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_C_XOR;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_D;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_D1;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_D2;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_D3;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_D4;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_D5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_D6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_DO5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_DO6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_D_CY;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X68Y80_D_XOR;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_A;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_A1;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_A2;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_A3;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_A4;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_A5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_A5Q;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_A6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_AMUX;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_AO5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_AO6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_AQ;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_AX;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_A_CY;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_A_XOR;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_B;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_B1;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_B2;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_B3;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_B4;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_B5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_B5Q;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_B6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_BMUX;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_BO5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_BO6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_BQ;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_BX;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_B_CY;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_B_XOR;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_C;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_C1;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_C2;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_C3;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_C4;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_C5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_C5Q;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_C6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_CE;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_CLK;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_CMUX;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_CO5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_CO6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_CQ;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_CX;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_C_CY;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_C_XOR;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_D;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_D1;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_D2;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_D3;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_D4;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_D5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_D5Q;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_D6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_DMUX;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_DO5;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_DO6;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_DQ;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_DX;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_D_CY;
  wire [0:0] CLBLL_L_X42Y80_SLICE_X69Y80_D_XOR;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_A;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_A1;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_A2;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_A3;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_A4;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_A5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_A6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_AO5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_AO6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_AQ;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_AX;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_A_CY;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_A_XOR;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_B;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_B1;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_B2;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_B3;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_B4;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_B5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_B6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_BMUX;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_BO5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_BO6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_BQ;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_BX;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_B_CY;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_B_XOR;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_C;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_C1;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_C2;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_C3;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_C4;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_C5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_C6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_CLK;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_CMUX;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_CO5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_CO6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_COUT;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_CX;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_C_CY;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_C_XOR;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_D;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_D1;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_D2;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_D3;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_D4;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_D5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_D6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_DMUX;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_DO5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_DO6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_DQ;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_DX;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_D_CY;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X68Y90_D_XOR;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_A;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_A1;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_A2;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_A3;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_A4;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_A5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_A6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_AMUX;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_AO5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_AO6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_A_CY;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_A_XOR;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_B;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_B1;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_B2;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_B3;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_B4;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_B5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_B6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_BMUX;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_BO5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_BO6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_B_CY;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_B_XOR;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_C;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_C1;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_C2;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_C3;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_C4;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_C5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_C6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_CE;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_CLK;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_CMUX;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_CO5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_CO6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_CQ;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_CX;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_C_CY;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_C_XOR;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_D;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_D1;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_D2;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_D3;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_D4;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_D5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_D6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_DMUX;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_DO5;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_DO6;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_D_CY;
  wire [0:0] CLBLL_L_X42Y90_SLICE_X69Y90_D_XOR;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_A;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_A1;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_A2;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_A3;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_A4;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_A5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_A6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_AMUX;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_AO5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_AO6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_AQ;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_AX;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_A_CY;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_A_XOR;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_B;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_B1;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_B2;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_B3;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_B4;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_B5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_B6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_BMUX;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_BO5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_BO6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_BQ;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_BX;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_B_CY;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_B_XOR;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_C;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_C1;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_C2;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_C3;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_C4;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_C5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_C6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_CIN;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_CLK;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_CMUX;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_CO5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_CO6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_COUT;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_CQ;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_CX;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_C_CY;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_C_XOR;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_D;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_D1;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_D2;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_D3;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_D4;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_D5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_D6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_DMUX;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_DO5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_DO6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_DQ;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_DX;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X68Y91_D_XOR;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_A;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_A1;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_A2;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_A3;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_A4;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_A5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_A6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_AMUX;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_AO5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_AO6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_AQ;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_AX;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_A_CY;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_A_XOR;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_B;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_B1;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_B2;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_B3;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_B4;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_B5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_B6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_BO5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_BO6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_BQ;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_B_CY;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_B_XOR;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_C;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_C1;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_C2;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_C3;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_C4;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_C5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_C6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_CLK;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_CO5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_CO6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_CQ;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_C_CY;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_C_XOR;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_D;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_D1;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_D2;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_D3;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_D4;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_D5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_D5Q;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_D6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_DMUX;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_DO5;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_DO6;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_DQ;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_DX;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_D_CY;
  wire [0:0] CLBLL_L_X42Y91_SLICE_X69Y91_D_XOR;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_A;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_A1;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_A2;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_A3;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_A4;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_A5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_A6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_AMUX;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_AO5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_AO6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_AQ;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_AX;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_A_CY;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_A_XOR;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_B;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_B1;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_B2;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_B3;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_B4;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_B5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_B6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_BMUX;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_BO5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_BO6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_BQ;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_BX;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_B_CY;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_B_XOR;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_C;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_C1;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_C2;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_C3;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_C4;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_C5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_C6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_CE;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_CIN;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_CLK;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_CMUX;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_CO5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_CO6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_COUT;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_CQ;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_CX;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_C_CY;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_C_XOR;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_D;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_D1;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_D2;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_D3;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_D4;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_D5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_D5Q;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_D6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_DMUX;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_DO5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_DO6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_DX;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X68Y92_D_XOR;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_A;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_A1;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_A2;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_A3;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_A4;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_A5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_A6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_AMUX;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_AO5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_AO6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_AQ;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_A_CY;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_A_XOR;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_B;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_B1;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_B2;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_B3;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_B4;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_B5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_B5Q;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_B6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_BMUX;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_BO5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_BO6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_BQ;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_BX;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_B_CY;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_B_XOR;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_C;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_C1;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_C2;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_C3;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_C4;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_C5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_C5Q;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_C6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_CLK;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_CMUX;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_CO5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_CO6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_C_CY;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_C_XOR;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_D;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_D1;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_D2;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_D3;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_D4;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_D5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_D6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_DO5;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_DO6;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_DQ;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_D_CY;
  wire [0:0] CLBLL_L_X42Y92_SLICE_X69Y92_D_XOR;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_A;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_A1;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_A2;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_A3;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_A4;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_A5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_A5Q;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_A6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_AMUX;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_AO5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_AO6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_AX;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_A_CY;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_A_XOR;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_B;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_B1;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_B2;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_B3;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_B4;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_B5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_B6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_BMUX;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_BO5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_BO6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_BQ;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_BX;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_B_CY;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_B_XOR;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_C;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_C1;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_C2;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_C3;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_C4;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_C5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_C6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_CE;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_CLK;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_CMUX;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_CO5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_CO6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_COUT;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_CQ;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_CX;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_C_CY;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_C_XOR;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_D;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_D1;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_D2;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_D3;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_D4;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_D5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_D6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_DMUX;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_DO5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_DO6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_DQ;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_DX;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_D_CY;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_D_XOR;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X68Y93_SR;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_A;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_A1;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_A2;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_A3;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_A4;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_A5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_A6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_AMUX;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_AO5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_AO6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_A_CY;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_A_XOR;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_B;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_B1;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_B2;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_B3;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_B4;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_B5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_B6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_BMUX;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_BO5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_BO6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_BQ;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_BX;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_B_CY;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_B_XOR;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_C;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_C1;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_C2;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_C3;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_C4;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_C5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_C6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_CLK;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_CMUX;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_CO5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_CO6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_C_CY;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_C_XOR;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_D;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_D1;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_D2;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_D3;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_D4;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_D5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_D6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_DMUX;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_DO5;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_DO6;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_D_CY;
  wire [0:0] CLBLL_L_X42Y93_SLICE_X69Y93_D_XOR;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_A;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_A1;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_A2;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_A3;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_A4;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_A5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_A6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_AMUX;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_AO5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_AO6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_AX;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_A_CY;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_A_XOR;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_B;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_B1;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_B2;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_B3;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_B4;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_B5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_B6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_BMUX;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_BO5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_BO6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_BQ;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_BX;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_B_CY;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_B_XOR;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_C;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_C1;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_C2;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_C3;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_C4;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_C5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_C6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_CIN;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_CLK;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_CMUX;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_CO5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_CO6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_COUT;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_CX;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_C_CY;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_C_XOR;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_D;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_D1;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_D2;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_D3;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_D4;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_D5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_D6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_DMUX;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_DO5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_DO6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_DX;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X68Y94_D_XOR;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_A;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_A1;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_A2;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_A3;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_A4;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_A5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_A6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_AMUX;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_AO5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_AO6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_A_CY;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_A_XOR;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_B;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_B1;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_B2;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_B3;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_B4;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_B5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_B6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_BMUX;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_BO5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_BO6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_B_CY;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_B_XOR;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_C;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_C1;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_C2;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_C3;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_C4;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_C5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_C6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_CLK;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_CO5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_CO6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_CX;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_C_CY;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_C_XOR;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_D;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_D1;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_D2;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_D3;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_D4;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_D5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_D6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_DMUX;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_DO5;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_DO6;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_D_CY;
  wire [0:0] CLBLL_L_X42Y94_SLICE_X69Y94_D_XOR;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_A;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_A1;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_A2;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_A3;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_A4;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_A5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_A6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_AMUX;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_AO5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_AO6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_AX;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_A_CY;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_A_XOR;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_B;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_B1;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_B2;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_B3;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_B4;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_B5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_B6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_BMUX;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_BO5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_BO6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_BX;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_B_CY;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_B_XOR;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_C;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_C1;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_C2;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_C3;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_C4;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_C5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_C6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_CIN;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_CLK;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_CMUX;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_CO5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_CO6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_COUT;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_CX;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_C_CY;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_C_XOR;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_D;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_D1;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_D2;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_D3;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_D4;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_D5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_D5Q;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_D6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_DMUX;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_DO5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_DO6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_DX;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X68Y95_D_XOR;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_A;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_A1;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_A2;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_A3;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_A4;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_A5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_A5Q;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_A6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_AMUX;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_AO5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_AO6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_AQ;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_AX;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_A_CY;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_A_XOR;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_B;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_B1;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_B2;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_B3;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_B4;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_B5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_B6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_BO5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_BO6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_BQ;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_B_CY;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_B_XOR;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_C;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_C1;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_C2;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_C3;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_C4;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_C5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_C6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_CLK;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_CMUX;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_CO5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_CO6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_CQ;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_C_CY;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_C_XOR;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_D;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_D1;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_D2;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_D3;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_D4;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_D5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_D5Q;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_D6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_DMUX;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_DO5;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_DO6;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_DQ;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_DX;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_D_CY;
  wire [0:0] CLBLL_L_X42Y95_SLICE_X69Y95_D_XOR;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_A;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_A1;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_A2;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_A3;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_A4;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_A5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_A6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_AMUX;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_AO5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_AO6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_AQ;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_AX;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_A_CY;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_A_XOR;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_B;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_B1;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_B2;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_B3;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_B4;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_B5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_B6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_BMUX;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_BO5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_BQ;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_BX;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_B_CY;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_B_XOR;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_C;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_C1;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_C2;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_C3;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_C4;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_C5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_C6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_CLK;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_CMUX;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_CO5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_CO6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_CQ;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_CX;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_C_CY;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_C_XOR;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_D;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_D1;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_D2;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_D3;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_D4;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_D5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_D6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_DMUX;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_DO5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_DO6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_DQ;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_DX;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_D_CY;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X68Y96_D_XOR;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_A;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_A1;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_A2;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_A3;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_A4;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_A5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_A6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_AMUX;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_AO5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_AO6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_A_CY;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_A_XOR;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_B;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_B1;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_B2;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_B3;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_B4;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_B5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_B5Q;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_B6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_BMUX;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_BO5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_BQ;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_BX;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_B_CY;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_B_XOR;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_C;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_C1;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_C2;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_C3;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_C4;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_C5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_C6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_CLK;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_CMUX;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_CO5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_CO6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_C_CY;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_C_XOR;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_D;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_D1;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_D2;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_D3;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_D4;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_D5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_D6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_DMUX;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_DO5;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_DO6;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_D_CY;
  wire [0:0] CLBLL_L_X42Y96_SLICE_X69Y96_D_XOR;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_A;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_A1;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_A2;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_A3;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_A4;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_A5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_A6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_AMUX;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_AO5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_AO6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_AQ;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_A_CY;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_A_XOR;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_B;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_B1;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_B2;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_B3;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_B4;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_B5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_B6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_BMUX;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_BO5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_BO6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_BQ;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_BX;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_B_CY;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_B_XOR;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_C;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_C1;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_C2;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_C3;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_C4;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_C5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_C6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_CLK;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_CMUX;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_CO5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_C_CY;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_C_XOR;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_D;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_D1;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_D2;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_D3;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_D4;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_D5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_D6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_DMUX;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_DO5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_DO6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_D_CY;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X68Y97_D_XOR;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_A;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_A1;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_A2;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_A3;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_A4;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_A5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_A6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_AMUX;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_AO5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_AO6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_A_CY;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_A_XOR;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_B;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_B1;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_B2;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_B3;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_B4;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_B5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_B6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_BMUX;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_BO5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_BO6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_B_CY;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_B_XOR;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_C;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_C1;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_C2;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_C3;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_C4;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_C5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_C5Q;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_C6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_CE;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_CLK;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_CMUX;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_CO5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_CO6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_C_CY;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_C_XOR;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_D;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_D1;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_D2;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_D3;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_D4;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_D5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_D6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_DMUX;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_DO5;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_DO6;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_D_CY;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_D_XOR;
  wire [0:0] CLBLL_L_X42Y97_SLICE_X69Y97_SR;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_A;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_A1;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_A2;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_A3;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_A4;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_A5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_A6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_AO5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_AO6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_A_CY;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_A_XOR;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_B;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_B1;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_B2;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_B3;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_B4;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_B5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_B6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_BO5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_BO6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_B_CY;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_B_XOR;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_C;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_C1;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_C2;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_C3;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_C4;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_C5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_C6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_CO5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_CO6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_C_CY;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_C_XOR;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_D;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_D1;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_D2;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_D3;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_D4;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_D5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_D6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_DO5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_DO6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_D_CY;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X68Y98_D_XOR;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_A;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_A1;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_A2;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_A3;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_A4;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_A5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_A6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_AO5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_AO6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_A_CY;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_A_XOR;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_B;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_B1;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_B2;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_B3;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_B4;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_B5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_B6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_BO5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_BO6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_BQ;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_BX;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_B_CY;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_B_XOR;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_C;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_C1;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_C2;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_C3;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_C4;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_C5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_C6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_CE;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_CLK;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_CO5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_CO6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_C_CY;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_C_XOR;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_D;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_D1;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_D2;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_D3;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_D4;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_D5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_D5Q;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_D6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_DMUX;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_DO5;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_DO6;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_DX;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_D_CY;
  wire [0:0] CLBLL_L_X42Y98_SLICE_X69Y98_D_XOR;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_A;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_A1;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_A2;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_A3;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_A4;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_A5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_A6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_AO5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_AO6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_A_CY;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_A_XOR;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_B;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_B1;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_B2;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_B3;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_B4;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_B5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_B6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_BO5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_BO6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_B_CY;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_B_XOR;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_C;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_C1;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_C2;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_C3;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_C4;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_C5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_C6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_CO5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_CO6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_C_CY;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_C_XOR;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_D;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_D1;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_D2;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_D3;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_D4;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_D5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_D6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_DO5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_DO6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_D_CY;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X2Y54_D_XOR;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_A;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_A1;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_A2;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_A3;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_A4;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_A5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_A6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_AMUX;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_AO5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_AO6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_AX;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_A_CY;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_A_XOR;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_B;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_B1;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_B2;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_B3;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_B4;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_B5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_B5Q;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_B6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_BMUX;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_BO5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_BO6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_BQ;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_BX;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_B_CY;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_B_XOR;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_C;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_C1;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_C2;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_C3;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_C4;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_C5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_C6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_CLK;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_CO5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_CO6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_COUT;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_CQ;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_CX;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_C_CY;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_C_XOR;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_D;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_D1;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_D2;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_D3;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_D4;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_D5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_D6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_DO5;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_DO6;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_DQ;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_DX;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_D_CY;
  wire [0:0] CLBLM_R_X3Y54_SLICE_X3Y54_D_XOR;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_A;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_A1;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_A2;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_A3;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_A4;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_A5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_A6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_AO5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_AO6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_A_CY;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_A_XOR;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_B;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_B1;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_B2;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_B3;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_B4;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_B5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_B6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_BO5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_BO6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_B_CY;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_B_XOR;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_C;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_C1;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_C2;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_C3;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_C4;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_C5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_C6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_CO5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_CO6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_C_CY;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_C_XOR;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_D;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_D1;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_D2;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_D3;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_D4;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_D5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_D6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_DO5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_DO6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_D_CY;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X2Y55_D_XOR;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_A;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_A1;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_A2;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_A3;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_A4;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_A5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_A6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_AMUX;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_AO5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_AO6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_AQ;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_AX;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_A_CY;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_A_XOR;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_B;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_B1;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_B2;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_B3;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_B4;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_B5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_B5Q;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_B6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_BMUX;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_BO5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_BO6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_BQ;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_BX;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_B_CY;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_B_XOR;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_C;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_C1;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_C2;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_C3;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_C4;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_C5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_C6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_CIN;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_CLK;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_CMUX;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_CO5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_CO6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_COUT;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_CX;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_C_CY;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_C_XOR;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_D;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_D1;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_D2;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_D3;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_D4;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_D5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_D6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_DMUX;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_DO5;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_DO6;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_DQ;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_DX;
  wire [0:0] CLBLM_R_X3Y55_SLICE_X3Y55_D_XOR;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_A;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_A1;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_A2;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_A3;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_A4;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_A5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_A6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_AO5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_AO6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_A_CY;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_A_XOR;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_B;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_B1;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_B2;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_B3;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_B4;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_B5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_B6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_BO5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_BO6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_B_CY;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_B_XOR;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_C;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_C1;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_C2;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_C3;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_C4;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_C5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_C6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_CO5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_CO6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_C_CY;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_C_XOR;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_D;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_D1;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_D2;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_D3;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_D4;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_D5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_D6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_DO5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_DO6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_D_CY;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X2Y56_D_XOR;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_A;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_A1;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_A2;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_A3;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_A4;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_A5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_A6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_AMUX;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_AO5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_AO6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_AQ;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_AX;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_A_CY;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_A_XOR;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_B;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_B1;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_B2;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_B3;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_B4;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_B5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_B5Q;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_B6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_BMUX;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_BO5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_BO6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_BQ;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_BX;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_B_CY;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_B_XOR;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_C;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_C1;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_C2;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_C3;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_C4;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_C5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_C6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_CIN;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_CLK;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_CMUX;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_CO5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_CO6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_COUT;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_CX;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_C_CY;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_C_XOR;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_D;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_D1;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_D2;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_D3;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_D4;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_D5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_D6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_DMUX;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_DO5;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_DO6;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_DQ;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_DX;
  wire [0:0] CLBLM_R_X3Y56_SLICE_X3Y56_D_XOR;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_A;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_A1;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_A2;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_A3;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_A4;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_A5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_A6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_AO5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_AO6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_A_CY;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_A_XOR;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_B;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_B1;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_B2;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_B3;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_B4;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_B5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_B6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_BO5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_BO6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_B_CY;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_B_XOR;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_C;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_C1;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_C2;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_C3;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_C4;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_C5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_C6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_CO5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_CO6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_C_CY;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_C_XOR;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_D;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_D1;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_D2;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_D3;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_D4;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_D5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_D6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_DO5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_DO6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_D_CY;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X2Y57_D_XOR;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_A;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_A1;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_A2;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_A3;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_A4;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_A5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_A6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_AMUX;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_AO5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_AO6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_AQ;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_AX;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_A_CY;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_A_XOR;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_B;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_B1;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_B2;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_B3;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_B4;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_B5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_B5Q;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_B6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_BMUX;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_BO5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_BO6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_BQ;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_BX;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_B_CY;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_B_XOR;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_C;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_C1;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_C2;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_C3;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_C4;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_C5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_C6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_CIN;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_CLK;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_CMUX;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_CO5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_CO6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_COUT;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_CX;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_C_CY;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_C_XOR;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_D;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_D1;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_D2;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_D3;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_D4;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_D5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_D6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_DMUX;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_DO5;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_DO6;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_DQ;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_DX;
  wire [0:0] CLBLM_R_X3Y57_SLICE_X3Y57_D_XOR;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_A;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_A1;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_A2;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_A3;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_A4;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_A5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_A6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_AO5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_AO6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_A_CY;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_A_XOR;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_B;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_B1;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_B2;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_B3;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_B4;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_B5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_B6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_BO5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_BO6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_B_CY;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_B_XOR;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_C;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_C1;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_C2;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_C3;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_C4;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_C5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_C6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_CO5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_CO6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_C_CY;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_C_XOR;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_D;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_D1;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_D2;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_D3;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_D4;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_D5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_D6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_DO5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_DO6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_D_CY;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X2Y58_D_XOR;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_A;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_A1;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_A2;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_A3;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_A4;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_A5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_A6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_AMUX;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_AO5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_AO6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_AQ;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_AX;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_A_CY;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_A_XOR;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_B;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_B1;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_B2;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_B3;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_B4;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_B5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_B5Q;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_B6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_BMUX;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_BO5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_BO6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_BQ;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_BX;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_B_CY;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_B_XOR;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_C;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_C1;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_C2;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_C3;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_C4;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_C5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_C6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_CIN;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_CLK;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_CMUX;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_CO5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_CO6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_COUT;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_CX;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_C_CY;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_C_XOR;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_D;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_D1;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_D2;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_D3;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_D4;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_D5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_D6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_DMUX;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_DO5;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_DO6;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_DQ;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_DX;
  wire [0:0] CLBLM_R_X3Y58_SLICE_X3Y58_D_XOR;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_A;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_A1;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_A2;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_A3;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_A4;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_A5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_A6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_AO5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_AO6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_A_CY;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_A_XOR;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_B;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_B1;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_B2;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_B3;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_B4;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_B5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_B6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_BO5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_BO6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_B_CY;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_B_XOR;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_C;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_C1;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_C2;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_C3;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_C4;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_C5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_C6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_CO5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_CO6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_C_CY;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_C_XOR;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_D;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_D1;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_D2;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_D3;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_D4;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_D5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_D6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_DO5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_DO6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_D_CY;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X2Y59_D_XOR;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_A;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_A1;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_A2;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_A3;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_A4;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_A5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_A6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_AMUX;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_AO5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_AO6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_AQ;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_AX;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_A_CY;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_A_XOR;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_B;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_B1;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_B2;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_B3;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_B4;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_B5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_B5Q;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_B6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_BMUX;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_BO5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_BO6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_BQ;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_BX;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_B_CY;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_B_XOR;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_C;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_C1;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_C2;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_C3;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_C4;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_C5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_C6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_CIN;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_CLK;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_CMUX;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_CO5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_CO6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_COUT;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_CX;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_C_CY;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_C_XOR;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_D;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_D1;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_D2;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_D3;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_D4;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_D5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_D6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_DMUX;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_DO5;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_DO6;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_DQ;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_DX;
  wire [0:0] CLBLM_R_X3Y59_SLICE_X3Y59_D_XOR;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_A;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_A1;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_A2;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_A3;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_A4;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_A5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_A6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_AO5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_AO6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_A_CY;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_A_XOR;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_B;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_B1;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_B2;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_B3;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_B4;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_B5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_B6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_BO5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_BO6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_B_CY;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_B_XOR;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_C;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_C1;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_C2;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_C3;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_C4;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_C5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_C6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_CO5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_CO6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_C_CY;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_C_XOR;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_D;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_D1;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_D2;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_D3;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_D4;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_D5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_D6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_DO5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_DO6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_D_CY;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X2Y60_D_XOR;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_A;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_A1;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_A2;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_A3;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_A4;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_A5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_A6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_AMUX;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_AO5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_AO6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_AX;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_A_CY;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_A_XOR;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_B;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_B1;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_B2;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_B3;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_B4;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_B5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_B5Q;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_B6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_BMUX;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_BO5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_BO6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_BQ;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_BX;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_B_CY;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_B_XOR;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_C;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_C1;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_C2;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_C3;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_C4;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_C5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_C6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_CIN;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_CLK;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_CO5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_CO6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_COUT;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_CX;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_C_CY;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_C_XOR;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_D;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_D1;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_D2;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_D3;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_D4;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_D5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_D6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_DO5;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_DO6;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_DX;
  wire [0:0] CLBLM_R_X3Y60_SLICE_X3Y60_D_XOR;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_A;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_A1;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_A2;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_A3;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_A4;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_A5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_A6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_AO5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_AO6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_A_CY;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_A_XOR;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_B;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_B1;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_B2;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_B3;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_B4;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_B5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_B6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_BO5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_BO6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_B_CY;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_B_XOR;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_C;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_C1;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_C2;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_C3;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_C4;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_C5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_C6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_CO5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_CO6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_C_CY;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_C_XOR;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_D;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_D1;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_D2;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_D3;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_D4;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_D5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_D6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_DO5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_DO6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_D_CY;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X66Y100_D_XOR;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_A;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_A1;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_A2;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_A3;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_A4;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_A5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_A5Q;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_A6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_AMUX;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_AO5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_AO6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_AQ;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_AX;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_A_CY;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_A_XOR;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_B;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_B1;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_B2;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_B3;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_B4;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_B5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_B6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_BMUX;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_BO5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_BO6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_BQ;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_BX;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_B_CY;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_B_XOR;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_C;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_C1;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_C2;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_C3;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_C4;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_C5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_C5Q;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_C6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_CE;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_CLK;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_CMUX;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_CO5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_CO6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_CQ;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_CX;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_C_CY;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_C_XOR;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_D;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_D1;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_D2;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_D3;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_D4;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_D5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_D5Q;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_D6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_DMUX;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_DO5;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_DO6;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_DQ;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_DX;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_D_CY;
  wire [0:0] CLBLM_R_X41Y100_SLICE_X67Y100_D_XOR;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_A;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_A1;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_A2;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_A3;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_A4;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_A5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_A6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_AO5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_AO6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_A_CY;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_A_XOR;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_B;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_B1;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_B2;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_B3;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_B4;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_B5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_B6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_BMUX;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_BO5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_BO6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_B_CY;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_B_XOR;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_C;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_C1;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_C2;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_C3;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_C4;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_C5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_C6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_CMUX;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_CO5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_CO6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_C_CY;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_C_XOR;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_D;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_D1;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_D2;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_D3;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_D4;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_D5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_D6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_DMUX;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_DO5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_DO6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_D_CY;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X66Y101_D_XOR;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_A;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_A1;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_A2;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_A3;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_A4;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_A5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_A6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_AMUX;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_AO5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_AO6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_A_CY;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_A_XOR;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_B;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_B1;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_B2;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_B3;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_B4;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_B5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_B6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_BMUX;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_BO5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_BO6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_B_CY;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_B_XOR;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_C;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_C1;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_C2;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_C3;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_C4;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_C5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_C6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_CE;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_CLK;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_CMUX;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_CO5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_CO6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_CX;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_C_CY;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_C_XOR;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_D;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_D1;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_D2;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_D3;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_D4;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_D5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_D6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_DMUX;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_DO5;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_DO6;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_DX;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_D_CY;
  wire [0:0] CLBLM_R_X41Y101_SLICE_X67Y101_D_XOR;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_A;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_A1;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_A2;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_A3;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_A4;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_A5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_A6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_AMUX;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_AO5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_AO6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_A_CY;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_A_XOR;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_B;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_B1;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_B2;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_B3;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_B4;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_B5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_B6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_BMUX;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_BO5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_BO6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_BQ;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_BX;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_B_CY;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_B_XOR;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_C;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_C1;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_C2;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_C3;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_C4;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_C5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_C6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_CLK;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_CMUX;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_CO5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_CO6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_C_CY;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_C_XOR;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_D;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_D1;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_D2;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_D3;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_D4;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_D5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_D6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_DMUX;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_DO5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_DO6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_D_CY;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X66Y102_D_XOR;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_A;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_A1;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_A2;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_A3;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_A4;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_A5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_A6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_AMUX;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_AO5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_AO6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_A_CY;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_A_XOR;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_B;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_B1;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_B2;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_B3;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_B4;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_B5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_B6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_BMUX;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_BO5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_BO6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_B_CY;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_B_XOR;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_C;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_C1;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_C2;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_C3;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_C4;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_C5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_C5Q;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_C6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_CE;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_CLK;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_CMUX;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_CO5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_CO6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_C_CY;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_C_XOR;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_D;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_D1;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_D2;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_D3;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_D4;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_D5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_D6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_DMUX;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_DO5;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_DO6;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_D_CY;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_D_XOR;
  wire [0:0] CLBLM_R_X41Y102_SLICE_X67Y102_SR;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_A;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_A1;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_A2;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_A3;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_A4;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_A5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_A6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_AO5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_AO6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_A_CY;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_A_XOR;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_B;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_B1;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_B2;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_B3;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_B4;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_B5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_B6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_BMUX;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_BO5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_BO6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_B_CY;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_B_XOR;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_C;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_C1;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_C2;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_C3;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_C4;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_C5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_C6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_CMUX;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_CO5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_CO6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_C_CY;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_C_XOR;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_D;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_D1;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_D2;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_D3;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_D4;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_D5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_D6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_DO5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_DO6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_D_CY;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X66Y103_D_XOR;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_A;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_A1;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_A2;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_A3;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_A4;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_A5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_A6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_AMUX;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_AO5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_AO6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_A_CY;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_A_XOR;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_B;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_B1;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_B2;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_B3;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_B4;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_B5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_B6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_BMUX;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_BO5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_BO6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_B_CY;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_B_XOR;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_C;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_C1;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_C2;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_C3;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_C4;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_C5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_C6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_CE;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_CLK;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_CMUX;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_CO5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_CO6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_C_CY;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_C_XOR;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_D;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_D1;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_D2;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_D3;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_D4;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_D5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_D5Q;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_D6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_DMUX;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_DO5;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_DO6;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_D_CY;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_D_XOR;
  wire [0:0] CLBLM_R_X41Y103_SLICE_X67Y103_SR;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_A;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_A1;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_A2;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_A3;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_A4;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_A5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_A6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_AMUX;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_AO5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_AO6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_A_CY;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_A_XOR;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_B;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_B1;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_B2;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_B3;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_B4;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_B5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_B6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_BMUX;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_BO5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_BO6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_B_CY;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_B_XOR;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_C;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_C1;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_C2;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_C3;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_C4;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_C5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_C6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_CE;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_CLK;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_CMUX;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_CO5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_CO6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_C_CY;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_C_XOR;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_D;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_D1;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_D2;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_D3;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_D4;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_D5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_D5Q;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_D6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_DMUX;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_DO5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_DO6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_DX;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_D_CY;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_D_XOR;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X66Y104_SR;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_A;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_A1;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_A2;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_A3;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_A4;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_A5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_A6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_AMUX;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_AO5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_AO6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_A_CY;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_A_XOR;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_B;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_B1;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_B2;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_B3;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_B4;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_B5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_B6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_BMUX;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_BO5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_BO6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_B_CY;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_B_XOR;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_C;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_C1;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_C2;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_C3;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_C4;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_C5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_C5Q;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_C6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_CE;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_CLK;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_CMUX;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_CO5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_CO6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_CX;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_C_CY;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_C_XOR;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_D;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_D1;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_D2;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_D3;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_D4;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_D5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_D6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_DMUX;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_DO5;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_DO6;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_D_CY;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_D_XOR;
  wire [0:0] CLBLM_R_X41Y104_SLICE_X67Y104_SR;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_A;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_A1;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_A2;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_A3;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_A4;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_A5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_A6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_AMUX;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_AO5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_AO6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_A_CY;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_A_XOR;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_B;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_B1;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_B2;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_B3;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_B4;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_B5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_B6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_BMUX;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_BO5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_BO6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_B_CY;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_B_XOR;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_C;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_C1;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_C2;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_C3;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_C4;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_C5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_C6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_CE;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_CLK;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_CMUX;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_CO5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_CO6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_C_CY;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_C_XOR;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_D;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_D1;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_D2;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_D3;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_D4;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_D5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_D6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_DO5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_DO6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_DQ;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_D_CY;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_D_XOR;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X66Y105_SR;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_A;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_A1;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_A2;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_A3;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_A4;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_A5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_A6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_AMUX;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_AO5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_AO6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_A_CY;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_A_XOR;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_B;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_B1;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_B2;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_B3;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_B4;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_B5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_B6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_BMUX;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_BO5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_BO6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_B_CY;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_B_XOR;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_C;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_C1;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_C2;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_C3;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_C4;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_C5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_C6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_CMUX;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_CO5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_CO6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_C_CY;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_C_XOR;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_D;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_D1;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_D2;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_D3;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_D4;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_D5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_D6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_DMUX;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_DO5;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_DO6;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_D_CY;
  wire [0:0] CLBLM_R_X41Y105_SLICE_X67Y105_D_XOR;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_A;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_A1;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_A2;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_A3;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_A4;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_A5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_A6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_AMUX;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_AO5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_AO6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_A_CY;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_A_XOR;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_B;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_B1;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_B2;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_B3;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_B4;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_B5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_B6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_BMUX;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_BO5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_BO6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_B_CY;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_B_XOR;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_C;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_C1;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_C2;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_C3;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_C4;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_C5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_C6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_CMUX;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_CO5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_CO6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_C_CY;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_C_XOR;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_D;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_D1;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_D2;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_D3;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_D4;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_D5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_D6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_DMUX;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_DO5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_DO6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_D_CY;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X66Y106_D_XOR;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_A;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_A1;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_A2;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_A3;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_A4;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_A5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_A5Q;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_A6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_AMUX;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_AO5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_AO6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_AQ;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_AX;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_A_CY;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_A_XOR;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_B;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_B1;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_B2;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_B3;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_B4;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_B5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_B6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_BMUX;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_BO5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_BO6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_BQ;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_BX;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_B_CY;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_B_XOR;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_C;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_C1;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_C2;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_C3;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_C4;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_C5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_C5Q;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_C6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_CE;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_CLK;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_CMUX;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_CO5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_CO6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_CQ;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_CX;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_C_CY;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_C_XOR;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_D;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_D1;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_D2;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_D3;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_D4;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_D5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_D6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_DMUX;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_DO5;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_DO6;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_D_CY;
  wire [0:0] CLBLM_R_X41Y106_SLICE_X67Y106_D_XOR;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_A;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_A1;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_A2;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_A3;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_A4;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_A5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_A6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_AMUX;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_AO5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_AO6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_A_CY;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_A_XOR;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_B;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_B1;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_B2;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_B3;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_B4;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_B5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_B6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_BMUX;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_BO5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_BO6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_B_CY;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_B_XOR;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_C;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_C1;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_C2;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_C3;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_C4;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_C5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_C6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_CMUX;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_CO5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_CO6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_C_CY;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_C_XOR;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_D;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_D1;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_D2;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_D3;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_D4;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_D5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_D6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_DMUX;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_DO5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_DO6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_D_CY;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X66Y107_D_XOR;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_A;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_A1;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_A2;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_A3;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_A4;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_A5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_A6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_AMUX;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_AO5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_AO6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_A_CY;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_A_XOR;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_B;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_B1;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_B2;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_B3;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_B4;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_B5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_B6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_BMUX;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_BO5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_BO6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_B_CY;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_B_XOR;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_C;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_C1;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_C2;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_C3;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_C4;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_C5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_C6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_CE;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_CLK;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_CMUX;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_CO5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_CO6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_C_CY;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_C_XOR;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_D;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_D1;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_D2;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_D3;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_D4;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_D5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_D5Q;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_D6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_DMUX;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_DO5;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_DO6;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_DX;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_D_CY;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_D_XOR;
  wire [0:0] CLBLM_R_X41Y107_SLICE_X67Y107_SR;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_A;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_A1;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_A2;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_A3;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_A4;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_A5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_A6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_AMUX;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_AO5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_AO6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_A_CY;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_A_XOR;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_B;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_B1;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_B2;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_B3;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_B4;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_B5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_B6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_BMUX;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_BO5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_BO6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_B_CY;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_B_XOR;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_C;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_C1;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_C2;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_C3;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_C4;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_C5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_C6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_CE;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_CLK;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_CMUX;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_CO5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_CO6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_C_CY;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_C_XOR;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_D;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_D1;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_D2;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_D3;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_D4;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_D5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_D5Q;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_D6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_DMUX;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_DO5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_DO6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_DX;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_D_CY;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_D_XOR;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X66Y108_SR;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_A;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_A1;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_A2;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_A3;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_A4;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_A5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_A6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_AMUX;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_AO5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_AO6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_A_CY;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_A_XOR;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_B;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_B1;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_B2;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_B3;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_B4;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_B5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_B6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_BMUX;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_BO5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_BO6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_B_CY;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_B_XOR;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_C;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_C1;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_C2;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_C3;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_C4;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_C5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_C6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_CLK;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_CMUX;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_CO5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_CO6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_C_CY;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_C_XOR;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_D;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_D1;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_D2;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_D3;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_D4;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_D5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_D5Q;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_D6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_DMUX;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_DO5;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_DO6;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_DX;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_D_CY;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_D_XOR;
  wire [0:0] CLBLM_R_X41Y108_SLICE_X67Y108_SR;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_A;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_A1;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_A2;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_A3;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_A4;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_A5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_A6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_AO5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_AO6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_AQ;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_A_CY;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_A_XOR;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_B;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_B1;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_B2;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_B3;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_B4;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_B5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_B6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_BMUX;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_BO5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_BO6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_B_CY;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_B_XOR;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_C;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_C1;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_C2;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_C3;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_C4;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_C5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_C6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_CE;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_CLK;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_CMUX;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_CO5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_CO6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_C_CY;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_C_XOR;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_D;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_D1;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_D2;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_D3;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_D4;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_D5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_D6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_DMUX;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_DO5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_DO6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_D_CY;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_D_XOR;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X66Y109_SR;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_A;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_A1;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_A2;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_A3;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_A4;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_A5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_A6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_AMUX;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_AO5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_AO6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_A_CY;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_A_XOR;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_B;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_B1;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_B2;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_B3;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_B4;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_B5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_B6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_BMUX;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_BO5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_BO6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_B_CY;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_B_XOR;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_C;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_C1;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_C2;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_C3;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_C4;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_C5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_C6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_CE;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_CLK;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_CMUX;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_CO5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_CO6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_C_CY;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_C_XOR;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_D;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_D1;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_D2;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_D3;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_D4;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_D5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_D5Q;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_D6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_DMUX;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_DO5;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_DO6;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_D_CY;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_D_XOR;
  wire [0:0] CLBLM_R_X41Y109_SLICE_X67Y109_SR;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_A;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_A1;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_A2;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_A3;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_A4;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_A5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_A6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_AMUX;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_AO5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_AO6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_A_CY;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_A_XOR;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_B;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_B1;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_B2;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_B3;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_B4;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_B5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_B5Q;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_B6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_BMUX;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_BO5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_BO6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_B_CY;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_B_XOR;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_C;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_C1;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_C2;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_C3;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_C4;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_C5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_C6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_CE;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_CLK;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_CMUX;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_CO5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_CO6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_C_CY;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_C_XOR;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_D;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_D1;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_D2;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_D3;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_D4;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_D5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_D6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_DMUX;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_DO5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_DO6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_D_CY;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_D_XOR;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X66Y110_SR;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_A;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_A1;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_A2;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_A3;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_A4;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_A5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_A6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_AMUX;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_AO5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_AO6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_A_CY;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_A_XOR;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_B;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_B1;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_B2;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_B3;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_B4;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_B5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_B5Q;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_B6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_BMUX;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_BO5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_BO6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_B_CY;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_B_XOR;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_C;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_C1;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_C2;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_C3;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_C4;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_C5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_C6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_CE;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_CLK;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_CMUX;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_CO5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_CO6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_C_CY;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_C_XOR;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_D;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_D1;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_D2;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_D3;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_D4;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_D5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_D6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_DMUX;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_DO5;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_DO6;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_D_CY;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_D_XOR;
  wire [0:0] CLBLM_R_X41Y110_SLICE_X67Y110_SR;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_A;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_A1;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_A2;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_A3;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_A4;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_A5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_A5Q;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_A6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_AMUX;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_AO5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_AO6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_AQ;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_AX;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_A_CY;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_A_XOR;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_B;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_B1;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_B2;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_B3;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_B4;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_B5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_B6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_BMUX;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_BO5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_BO6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_BQ;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_BX;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_B_CY;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_B_XOR;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_C;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_C1;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_C2;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_C3;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_C4;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_C5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_C6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_CE;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_CLK;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_CMUX;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_CO5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_CO6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_C_CY;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_C_XOR;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_D;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_D1;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_D2;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_D3;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_D4;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_D5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_D6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_DMUX;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_DO5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_DO6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_DQ;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_DX;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_D_CY;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X66Y111_D_XOR;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_A;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_A1;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_A2;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_A3;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_A4;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_A5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_A5Q;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_A6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_AMUX;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_AO5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_AO6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_A_CY;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_A_XOR;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_B;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_B1;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_B2;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_B3;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_B4;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_B5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_B6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_BMUX;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_BO5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_BO6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_B_CY;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_B_XOR;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_C;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_C1;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_C2;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_C3;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_C4;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_C5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_C6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_CE;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_CLK;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_CMUX;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_CO5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_CO6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_C_CY;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_C_XOR;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_D;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_D1;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_D2;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_D3;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_D4;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_D5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_D6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_DMUX;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_DO5;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_DO6;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_D_CY;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_D_XOR;
  wire [0:0] CLBLM_R_X41Y111_SLICE_X67Y111_SR;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_A;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_A1;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_A2;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_A3;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_A4;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_A5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_A6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_AMUX;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_AO5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_AO6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_A_CY;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_A_XOR;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_B;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_B1;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_B2;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_B3;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_B4;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_B5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_B6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_BMUX;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_BO5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_BO6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_B_CY;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_B_XOR;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_C;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_C1;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_C2;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_C3;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_C4;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_C5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_C6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_CLK;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_CO5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_CO6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_CQ;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_C_CY;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_C_XOR;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_D;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_D1;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_D2;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_D3;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_D4;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_D5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_D5Q;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_D6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_DMUX;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_DO5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_DO6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_DQ;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_DX;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_D_CY;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X66Y114_D_XOR;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_A;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_A1;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_A2;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_A3;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_A4;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_A5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_A5Q;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_A6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_AMUX;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_AO5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_AO6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_AX;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_A_CY;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_A_XOR;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_B;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_B1;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_B2;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_B3;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_B4;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_B5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_B5Q;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_B6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_BMUX;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_BO5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_BO6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_BX;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_B_CY;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_B_XOR;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_C;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_C1;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_C2;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_C3;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_C4;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_C5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_C6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_CE;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_CLK;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_CMUX;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_CO5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_CO6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_COUT;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_CQ;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_CX;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_C_CY;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_C_XOR;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_D;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_D1;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_D2;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_D3;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_D4;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_D5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_D6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_DMUX;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_DO5;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_DO6;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_DQ;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_DX;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_D_CY;
  wire [0:0] CLBLM_R_X41Y114_SLICE_X67Y114_D_XOR;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_A;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_A1;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_A2;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_A3;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_A4;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_A5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_A6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_AMUX;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_AO5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_AO6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_A_CY;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_A_XOR;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_B;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_B1;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_B2;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_B3;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_B4;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_B5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_B6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_BMUX;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_BO5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_BO6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_BQ;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_B_CY;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_B_XOR;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_C;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_C1;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_C2;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_C3;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_C4;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_C5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_C6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_CLK;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_CMUX;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_CO5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_CO6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_C_CY;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_C_XOR;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_D;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_D1;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_D2;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_D3;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_D4;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_D5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_D5Q;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_D6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_DMUX;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_DO5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_DO6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_DQ;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_DX;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_D_CY;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X66Y115_D_XOR;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_A;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_A1;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_A2;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_A3;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_A4;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_A5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_A6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_AMUX;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_AO5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_AO6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_AQ;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_AX;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_A_CY;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_A_XOR;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_B;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_B1;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_B2;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_B3;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_B4;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_B5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_B6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_BMUX;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_BO5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_BO6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_BQ;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_BX;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_B_CY;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_B_XOR;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_C;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_C1;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_C2;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_C3;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_C4;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_C5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_C6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_CE;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_CIN;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_CLK;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_CMUX;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_CO5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_CO6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_COUT;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_CQ;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_CX;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_C_CY;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_C_XOR;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_D;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_D1;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_D2;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_D3;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_D4;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_D5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_D6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_DMUX;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_DO5;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_DO6;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_DQ;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_DX;
  wire [0:0] CLBLM_R_X41Y115_SLICE_X67Y115_D_XOR;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_A;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_A1;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_A2;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_A3;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_A4;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_A5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_A6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_AMUX;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_AO5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_AO6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_A_CY;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_A_XOR;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_B;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_B1;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_B2;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_B3;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_B4;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_B5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_B6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_BMUX;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_BO5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_BO6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_B_CY;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_B_XOR;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_C;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_C1;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_C2;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_C3;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_C4;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_C5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_C6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_CLK;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_CO5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_CO6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_CQ;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_C_CY;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_C_XOR;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_D;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_D1;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_D2;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_D3;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_D4;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_D5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_D5Q;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_D6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_DMUX;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_DO5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_DO6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_DQ;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_DX;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_D_CY;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X66Y116_D_XOR;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_A;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_A1;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_A2;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_A3;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_A4;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_A5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_A6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_AMUX;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_AO5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_AO6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_AQ;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_AX;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_A_CY;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_B;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_B1;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_B2;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_B3;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_B4;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_B5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_B6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_BMUX;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_BO5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_BO6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_BX;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_B_CY;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_B_XOR;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_C;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_C1;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_C2;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_C3;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_C4;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_C5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_C6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_CE;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_CIN;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_CLK;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_CO5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_CO6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_COUT;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_CQ;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_CX;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_C_CY;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_C_XOR;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_D;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_D1;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_D2;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_D3;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_D4;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_D5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_D6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_DMUX;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_DO5;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_DO6;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_DX;
  wire [0:0] CLBLM_R_X41Y116_SLICE_X67Y116_D_XOR;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_A;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_A1;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_A2;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_A3;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_A4;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_A5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_A6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_AO5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_AO6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_A_CY;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_A_XOR;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_B;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_B1;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_B2;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_B3;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_B4;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_B5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_B6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_BO5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_BO6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_B_CY;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_B_XOR;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_C;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_C1;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_C2;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_C3;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_C4;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_C5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_C6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_CO5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_CO6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_C_CY;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_C_XOR;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_D;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_D1;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_D2;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_D3;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_D4;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_D5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_D6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_DO5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_DO6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_D_CY;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X66Y92_D_XOR;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_A;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_A1;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_A2;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_A3;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_A4;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_A5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_A6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_AMUX;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_AO5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_AO6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_AX;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_A_CY;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_A_XOR;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_B;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_B1;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_B2;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_B3;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_B4;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_B5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_B6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_BMUX;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_BO5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_BO6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_BQ;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_BX;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_B_CY;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_B_XOR;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_C;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_C1;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_C2;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_C3;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_C4;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_C5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_C6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_CE;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_CLK;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_CO5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_CO6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_COUT;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_CQ;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_CX;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_C_CY;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_C_XOR;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_D;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_D1;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_D2;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_D3;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_D4;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_D5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_D6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_DMUX;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_DO5;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_DO6;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_DQ;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_DX;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_D_CY;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_D_XOR;
  wire [0:0] CLBLM_R_X41Y92_SLICE_X67Y92_SR;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_A;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_A1;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_A2;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_A3;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_A4;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_A5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_A6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_AO5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_AO6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_A_CY;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_A_XOR;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_B;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_B1;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_B2;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_B3;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_B4;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_B5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_B6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_BO5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_BO6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_B_CY;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_B_XOR;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_C;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_C1;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_C2;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_C3;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_C4;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_C5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_C6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_CO5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_CO6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_C_CY;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_C_XOR;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_D;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_D1;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_D2;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_D3;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_D4;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_D5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_D6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_DO5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_DO6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_D_CY;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X66Y93_D_XOR;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_A;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_A1;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_A2;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_A3;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_A4;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_A5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_A5Q;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_A6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_AMUX;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_AO5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_AO6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_AQ;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_AX;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_A_CY;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_A_XOR;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_B;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_B1;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_B2;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_B3;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_B4;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_B5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_B5Q;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_B6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_BMUX;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_BO5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_BO6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_BQ;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_BX;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_B_CY;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_B_XOR;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_C;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_C1;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_C2;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_C3;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_C4;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_C5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_C5Q;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_C6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_CE;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_CIN;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_CLK;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_CMUX;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_CO5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_CO6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_COUT;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_CQ;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_CX;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_C_CY;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_C_XOR;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_D;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_D1;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_D2;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_D3;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_D4;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_D5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_D5Q;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_D6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_DMUX;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_DO5;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_DO6;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_DQ;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_DX;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_D_XOR;
  wire [0:0] CLBLM_R_X41Y93_SLICE_X67Y93_SR;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_A;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_A1;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_A2;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_A3;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_A4;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_A5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_A6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_AO5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_AO6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_A_CY;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_A_XOR;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_B;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_B1;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_B2;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_B3;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_B4;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_B5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_B6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_BO5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_BO6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_B_CY;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_B_XOR;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_C;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_C1;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_C2;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_C3;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_C4;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_C5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_C6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_CO5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_CO6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_C_CY;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_C_XOR;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_D;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_D1;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_D2;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_D3;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_D4;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_D5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_D6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_DO5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_DO6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_D_CY;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X66Y94_D_XOR;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_A;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_A1;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_A2;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_A3;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_A4;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_A5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_A6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_AMUX;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_AO5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_AO6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_AQ;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_AX;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_A_CY;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_A_XOR;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_B;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_B1;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_B2;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_B3;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_B4;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_B5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_B5Q;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_B6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_BMUX;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_BO5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_BO6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_BQ;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_BX;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_B_CY;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_B_XOR;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_C;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_C1;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_C2;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_C3;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_C4;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_C5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_C6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_CE;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_CIN;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_CLK;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_CMUX;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_CO5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_CO6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_COUT;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_CQ;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_CX;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_C_CY;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_C_XOR;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_D;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_D1;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_D2;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_D3;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_D4;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_D5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_D6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_DMUX;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_DO5;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_DO6;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_DQ;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_DX;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_D_XOR;
  wire [0:0] CLBLM_R_X41Y94_SLICE_X67Y94_SR;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_A;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_A1;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_A2;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_A3;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_A4;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_A5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_A6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_AO5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_AO6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_A_CY;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_A_XOR;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_B;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_B1;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_B2;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_B3;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_B4;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_B5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_B6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_BO5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_BO6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_B_CY;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_B_XOR;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_C;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_C1;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_C2;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_C3;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_C4;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_C5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_C6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_CO5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_CO6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_C_CY;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_C_XOR;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_D;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_D1;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_D2;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_D3;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_D4;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_D5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_D6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_DO5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_DO6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_D_CY;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X66Y95_D_XOR;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_A;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_A1;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_A2;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_A3;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_A4;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_A5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_A6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_AMUX;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_AO5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_AO6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_AQ;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_AX;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_A_CY;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_A_XOR;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_B;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_B1;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_B2;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_B3;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_B4;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_B5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_B6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_BMUX;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_BO5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_BO6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_BQ;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_BX;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_B_CY;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_B_XOR;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_C;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_C1;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_C2;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_C3;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_C4;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_C5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_C6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_CE;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_CIN;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_CLK;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_CMUX;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_CO5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_CO6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_COUT;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_CQ;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_CX;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_C_CY;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_C_XOR;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_D;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_D1;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_D2;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_D3;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_D4;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_D5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_D6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_DMUX;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_DO5;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_DO6;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_DQ;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_DX;
  wire [0:0] CLBLM_R_X41Y95_SLICE_X67Y95_D_XOR;
  wire [0:0] CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_CE0;
  wire [0:0] CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_CE1;
  wire [0:0] CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_I0;
  wire [0:0] CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_I1;
  wire [0:0] CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_IGNORE0;
  wire [0:0] CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_IGNORE1;
  wire [0:0] CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_O;
  wire [0:0] CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_S0;
  wire [0:0] CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_S1;
  wire [0:0] CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_CE;
  wire [0:0] CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_I;
  wire [0:0] CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O;
  wire [0:0] CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_CE;
  wire [0:0] CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_I;
  wire [0:0] CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  wire [0:0] CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_CE;
  wire [0:0] CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_I;
  wire [0:0] CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  wire [0:0] LIOB33_X0Y55_IOB_X0Y55_O;
  wire [0:0] LIOB33_X0Y57_IOB_X0Y57_O;
  wire [0:0] LIOB33_X0Y59_IOB_X0Y59_O;
  wire [0:0] LIOB33_X0Y67_IOB_X0Y68_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_TQ;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_D1;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_OQ;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_T1;
  wire [0:0] LIOI3_X0Y55_OLOGIC_X0Y55_TQ;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_D1;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_OQ;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_T1;
  wire [0:0] LIOI3_X0Y59_OLOGIC_X0Y59_TQ;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y68_D1;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y68_OQ;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y68_T1;
  wire [0:0] LIOI3_X0Y67_OLOGIC_X0Y68_TQ;
  wire [0:0] RIOB33_X57Y125_IOB_X1Y126_I;
  wire [0:0] RIOB33_X57Y127_IOB_X1Y127_O;
  wire [0:0] RIOI3_X57Y125_ILOGIC_X1Y126_D;
  wire [0:0] RIOI3_X57Y125_ILOGIC_X1Y126_O;
  wire [0:0] RIOI3_X57Y127_OLOGIC_X1Y127_D1;
  wire [0:0] RIOI3_X57Y127_OLOGIC_X1Y127_OQ;
  wire [0:0] RIOI3_X57Y127_OLOGIC_X1Y127_T1;
  wire [0:0] RIOI3_X57Y127_OLOGIC_X1Y127_TQ;


  (* KEEP, DONT_TOUCH, BEL = "RAMB18E1" *)
  RAMB18E1 #(
    .DOA_REG(0),
    .DOB_REG(0),
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h5555555555555555555555555555555555555555555555555555555555555555),
    .INITP_03(256'h5555555555555555555555555555555555555555555555555555555555555555),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h5555555555555555555555555555555555555555555555555555555555555555),
    .INITP_07(256'h5555555555555555555555555555555555555555555555555555555555555555),
    .INIT_00(256'h000F000E000D000C000B000A0009000800070006000500040003000200010000),
    .INIT_01(256'h001F001E001D001C001B001A0019001800170016001500140013001200110010),
    .INIT_02(256'h002F002E002D002C002B002A0029002800270026002500240023002200210020),
    .INIT_03(256'h003F003E003D003C003B003A0039003800370036003500340033003200310030),
    .INIT_04(256'h004F004E004D004C004B004A0049004800470046004500440043004200410040),
    .INIT_05(256'h005F005E005D005C005B005A0059005800570056005500540053005200510050),
    .INIT_06(256'h006F006E006D006C006B006A0069006800670066006500640063006200610060),
    .INIT_07(256'h007F007E007D007C007B007A0079007800770076007500740073007200710070),
    .INIT_08(256'h008F008E008D008C008B008A0089008800870086008500840083008200810080),
    .INIT_09(256'h009F009E009D009C009B009A0099009800970096009500940093009200910090),
    .INIT_0A(256'h00AF00AE00AD00AC00AB00AA00A900A800A700A600A500A400A300A200A100A0),
    .INIT_0B(256'h00BF00BE00BD00BC00BB00BA00B900B800B700B600B500B400B300B200B100B0),
    .INIT_0C(256'h00CF00CE00CD00CC00CB00CA00C900C800C700C600C500C400C300C200C100C0),
    .INIT_0D(256'h00DF00DE00DD00DC00DB00DA00D900D800D700D600D500D400D300D200D100D0),
    .INIT_0E(256'h00EF00EE00ED00EC00EB00EA00E900E800E700E600E500E400E300E200E100E0),
    .INIT_0F(256'h00FF00FE00FD00FC00FB00FA00F900F800F700F600F500F400F300F200F100F0),
    .INIT_10(256'h000F000E000D000C000B000A0009000800070006000500040003000200010000),
    .INIT_11(256'h001F001E001D001C001B001A0019001800170016001500140013001200110010),
    .INIT_12(256'h002F002E002D002C002B002A0029002800270026002500240023002200210020),
    .INIT_13(256'h003F003E003D003C003B003A0039003800370036003500340033003200310030),
    .INIT_14(256'h004F004E004D004C004B004A0049004800470046004500440043004200410040),
    .INIT_15(256'h005F005E005D005C005B005A0059005800570056005500540053005200510050),
    .INIT_16(256'h006F006E006D006C006B006A0069006800670066006500640063006200610060),
    .INIT_17(256'h007F007E007D007C007B007A0079007800770076007500740073007200710070),
    .INIT_18(256'h008F008E008D008C008B008A0089008800870086008500840083008200810080),
    .INIT_19(256'h009F009E009D009C009B009A0099009800970096009500940093009200910090),
    .INIT_1A(256'h00AF00AE00AD00AC00AB00AA00A900A800A700A600A500A400A300A200A100A0),
    .INIT_1B(256'h00BF00BE00BD00BC00BB00BA00B900B800B700B600B500B400B300B200B100B0),
    .INIT_1C(256'h00CF00CE00CD00CC00CB00CA00C900C800C700C600C500C400C300C200C100C0),
    .INIT_1D(256'h00DF00DE00DD00DC00DB00DA00D900D800D700D600D500D400D300D200D100D0),
    .INIT_1E(256'h00EF00EE00ED00EC00EB00EA00E900E800E700E600E500E400E300E200E100E0),
    .INIT_1F(256'h00FF00FE00FD00FC00FB00FA00F900F800F700F600F500F400F300F200F100F0),
    .INIT_20(256'h010F010E010D010C010B010A0109010801070106010501040103010201010100),
    .INIT_21(256'h011F011E011D011C011B011A0119011801170116011501140113011201110110),
    .INIT_22(256'h012F012E012D012C012B012A0129012801270126012501240123012201210120),
    .INIT_23(256'h013F013E013D013C013B013A0139013801370136013501340133013201310130),
    .INIT_24(256'h014F014E014D014C014B014A0149014801470146014501440143014201410140),
    .INIT_25(256'h015F015E015D015C015B015A0159015801570156015501540153015201510150),
    .INIT_26(256'h016F016E016D016C016B016A0169016801670166016501640163016201610160),
    .INIT_27(256'h017F017E017D017C017B017A0179017801770176017501740173017201710170),
    .INIT_28(256'h018F018E018D018C018B018A0189018801870186018501840183018201810180),
    .INIT_29(256'h019F019E019D019C019B019A0199019801970196019501940193019201910190),
    .INIT_2A(256'h01AF01AE01AD01AC01AB01AA01A901A801A701A601A501A401A301A201A101A0),
    .INIT_2B(256'h01BF01BE01BD01BC01BB01BA01B901B801B701B601B501B401B301B201B101B0),
    .INIT_2C(256'h01CF01CE01CD01CC01CB01CA01C901C801C701C601C501C401C301C201C101C0),
    .INIT_2D(256'h01DF01DE01DD01DC01DB01DA01D901D801D701D601D501D401D301D201D101D0),
    .INIT_2E(256'h01EF01EE01ED01EC01EB01EA01E901E801E701E601E501E401E301E201E101E0),
    .INIT_2F(256'h01FF01FE01FD01FC01FB01FA01F901F801F701F601F501F401F301F201F101F0),
    .INIT_30(256'h010F010E010D010C010B010A0109010801070106010501040103010201010100),
    .INIT_31(256'h011F011E011D011C011B011A0119011801170116011501140113011201110110),
    .INIT_32(256'h012F012E012D012C012B012A0129012801270126012501240123012201210120),
    .INIT_33(256'h013F013E013D013C013B013A0139013801370136013501340133013201310130),
    .INIT_34(256'h014F014E014D014C014B014A0149014801470146014501440143014201410140),
    .INIT_35(256'h015F015E015D015C015B015A0159015801570156015501540153015201510150),
    .INIT_36(256'h016F016E016D016C016B016A0169016801670166016501640163016201610160),
    .INIT_37(256'h017F017E017D017C017B017A0179017801770176017501740173017201710170),
    .INIT_38(256'h018F018E018D018C018B018A0189018801870186018501840183018201810180),
    .INIT_39(256'h019F019E019D019C019B019A0199019801970196019501940193019201910190),
    .INIT_3A(256'h01AF01AE01AD01AC01AB01AA01A901A801A701A601A501A401A301A201A101A0),
    .INIT_3B(256'h01BF01BE01BD01BC01BB01BA01B901B801B701B601B501B401B301B201B101B0),
    .INIT_3C(256'h01CF01CE01CD01CC01CB01CA01C901C801C701C601C501C401C301C201C101C0),
    .INIT_3D(256'h01DF01DE01DD01DC01DB01DA01D901D801D701D601D501D401D301D201D101D0),
    .INIT_3E(256'h01EF01EE01ED01EC01EB01EA01E901E801E701E601E501E401E301E201E101E0),
    .INIT_3F(256'h01FF01FE01FD01FC01FB01FA01F901F801F701F601F501F401F301F201F101F0),
    .INIT_A(18'h00000),
    .INIT_B(18'h00000),
    .IS_CLKARDCLK_INVERTED(0),
    .IS_CLKBWRCLK_INVERTED(1),
    .IS_ENARDEN_INVERTED(0),
    .IS_ENBWREN_INVERTED(0),
    .IS_RSTRAMARSTRAM_INVERTED(1),
    .IS_RSTRAMB_INVERTED(1),
    .IS_RSTREGARSTREG_INVERTED(1),
    .IS_RSTREGB_INVERTED(1),
    .RAM_MODE("TDP"),
    .READ_WIDTH_A(18),
    .READ_WIDTH_B(18),
    .SRVAL_A(18'h00000),
    .SRVAL_B(18'h00000),
    .WRITE_MODE_A("READ_FIRST"),
    .WRITE_MODE_B("READ_FIRST"),
    .WRITE_WIDTH_A(18),
    .WRITE_WIDTH_B(18)
  ) BRAM_L_X44Y95_RAMB18_X2Y38_RAMB18E1 (
.ADDRARDADDR({CLBLL_L_X42Y92_SLICE_X69Y92_DQ, CLBLL_L_X42Y92_SLICE_X69Y92_C5Q, CLBLL_L_X42Y91_SLICE_X68Y91_DQ, CLBLL_L_X42Y91_SLICE_X68Y91_CQ, CLBLL_L_X42Y91_SLICE_X68Y91_BQ, CLBLL_L_X42Y91_SLICE_X68Y91_AQ, CLBLL_L_X42Y90_SLICE_X68Y90_AQ, CLBLL_L_X42Y90_SLICE_X68Y90_DQ, CLBLL_L_X42Y90_SLICE_X68Y90_BQ, CLBLL_L_X42Y94_SLICE_X68Y94_BQ, 1'b0, 1'b0, 1'b0, 1'b0}),
.ADDRBWRADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CLKARDCLK(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CLKBWRCLK(1'b1),
.DIADI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.DIBDI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.DIPADIP({1'b0, 1'b0}),
.DIPBDIP({1'b0, 1'b0}),
.DOADO({BRAM_L_X44Y95_RAMB18_X2Y38_DO15, BRAM_L_X44Y95_RAMB18_X2Y38_DO14, BRAM_L_X44Y95_RAMB18_X2Y38_DO13, BRAM_L_X44Y95_RAMB18_X2Y38_DO12, BRAM_L_X44Y95_RAMB18_X2Y38_DO11, BRAM_L_X44Y95_RAMB18_X2Y38_DO10, BRAM_L_X44Y95_RAMB18_X2Y38_DO9, BRAM_L_X44Y95_RAMB18_X2Y38_DO8, BRAM_L_X44Y95_RAMB18_X2Y38_DO7, BRAM_L_X44Y95_RAMB18_X2Y38_DO6, BRAM_L_X44Y95_RAMB18_X2Y38_DO5, BRAM_L_X44Y95_RAMB18_X2Y38_DO4, BRAM_L_X44Y95_RAMB18_X2Y38_DO3, BRAM_L_X44Y95_RAMB18_X2Y38_DO2, BRAM_L_X44Y95_RAMB18_X2Y38_DO1, BRAM_L_X44Y95_RAMB18_X2Y38_DO0}),
.DOBDO({BRAM_L_X44Y95_RAMB18_X2Y38_DO31, BRAM_L_X44Y95_RAMB18_X2Y38_DO30, BRAM_L_X44Y95_RAMB18_X2Y38_DO29, BRAM_L_X44Y95_RAMB18_X2Y38_DO28, BRAM_L_X44Y95_RAMB18_X2Y38_DO27, BRAM_L_X44Y95_RAMB18_X2Y38_DO26, BRAM_L_X44Y95_RAMB18_X2Y38_DO25, BRAM_L_X44Y95_RAMB18_X2Y38_DO24, BRAM_L_X44Y95_RAMB18_X2Y38_DO23, BRAM_L_X44Y95_RAMB18_X2Y38_DO22, BRAM_L_X44Y95_RAMB18_X2Y38_DO21, BRAM_L_X44Y95_RAMB18_X2Y38_DO20, BRAM_L_X44Y95_RAMB18_X2Y38_DO19, BRAM_L_X44Y95_RAMB18_X2Y38_DO18, BRAM_L_X44Y95_RAMB18_X2Y38_DO17, BRAM_L_X44Y95_RAMB18_X2Y38_DO16}),
.DOPADOP({BRAM_L_X44Y95_RAMB18_X2Y38_DOP1, BRAM_L_X44Y95_RAMB18_X2Y38_DOP0}),
.DOPBDOP({BRAM_L_X44Y95_RAMB18_X2Y38_DOP3, BRAM_L_X44Y95_RAMB18_X2Y38_DOP2}),
.ENARDEN(1'b1),
.ENBWREN(1'b1),
.REGCEAREGCE(1'b1),
.REGCEB(1'b0),
.RSTRAMARSTRAM(1'b1),
.RSTRAMB(1'b1),
.RSTREGARSTREG(1'b1),
.RSTREGB(1'b1),
.WEA({1'b0, 1'b0}),
.WEBWE({1'b0, 1'b0})
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X42Y43_SLICE_X68Y43_CARRY4 (
.CI(1'b0),
.CO({CLBLL_L_X42Y43_SLICE_X68Y43_D_CY, CLBLL_L_X42Y43_SLICE_X68Y43_C_CY, CLBLL_L_X42Y43_SLICE_X68Y43_B_CY, CLBLL_L_X42Y43_SLICE_X68Y43_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({CLBLL_L_X42Y43_SLICE_X68Y43_D_XOR, CLBLL_L_X42Y43_SLICE_X68Y43_C_XOR, CLBLL_L_X42Y43_SLICE_X68Y43_B_XOR, CLBLL_L_X42Y43_SLICE_X68Y43_A_XOR}),
.S({CLBLL_L_X42Y43_SLICE_X68Y43_DO6, CLBLL_L_X42Y43_SLICE_X68Y43_CO6, CLBLL_L_X42Y43_SLICE_X68Y43_BO6, CLBLL_L_X42Y43_SLICE_X68Y43_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000000000)
  ) CLBLL_L_X42Y43_SLICE_X68Y43_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b0),
.I5(1'b1),
.O5(CLBLL_L_X42Y43_SLICE_X68Y43_DO5),
.O6(CLBLL_L_X42Y43_SLICE_X68Y43_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000000000)
  ) CLBLL_L_X42Y43_SLICE_X68Y43_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X42Y96_SLICE_X69Y96_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y43_SLICE_X68Y43_CO5),
.O6(CLBLL_L_X42Y43_SLICE_X68Y43_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLL_L_X42Y43_SLICE_X68Y43_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y96_SLICE_X69Y96_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y43_SLICE_X68Y43_BO5),
.O6(CLBLL_L_X42Y43_SLICE_X68Y43_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLL_L_X42Y43_SLICE_X68Y43_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y110_SLICE_X69Y110_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y43_SLICE_X68Y43_AO5),
.O6(CLBLL_L_X42Y43_SLICE_X68Y43_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y43_SLICE_X69Y43_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y43_SLICE_X69Y43_DO5),
.O6(CLBLL_L_X42Y43_SLICE_X69Y43_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y43_SLICE_X69Y43_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y43_SLICE_X69Y43_CO5),
.O6(CLBLL_L_X42Y43_SLICE_X69Y43_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y43_SLICE_X69Y43_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y43_SLICE_X69Y43_BO5),
.O6(CLBLL_L_X42Y43_SLICE_X69Y43_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y43_SLICE_X69Y43_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y43_SLICE_X69Y43_AO5),
.O6(CLBLL_L_X42Y43_SLICE_X69Y43_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y68_SLICE_X68Y68_A5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y68_SLICE_X68Y68_AO5),
.Q(CLBLL_L_X42Y68_SLICE_X68Y68_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y68_SLICE_X68Y68_B5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y68_SLICE_X68Y68_BO5),
.Q(CLBLL_L_X42Y68_SLICE_X68Y68_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y68_SLICE_X68Y68_C5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y68_SLICE_X68Y68_CO5),
.Q(CLBLL_L_X42Y68_SLICE_X68Y68_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y68_SLICE_X68Y68_D5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y68_SLICE_X68Y68_DO5),
.Q(CLBLL_L_X42Y68_SLICE_X68Y68_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y68_SLICE_X68Y68_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y80_SLICE_X69Y80_D5Q),
.Q(CLBLL_L_X42Y68_SLICE_X68Y68_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y68_SLICE_X68Y68_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y80_SLICE_X69Y80_C5Q),
.Q(CLBLL_L_X42Y68_SLICE_X68Y68_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y68_SLICE_X68Y68_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y80_SLICE_X69Y80_DQ),
.Q(CLBLL_L_X42Y68_SLICE_X68Y68_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y68_SLICE_X68Y68_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y80_SLICE_X69Y80_AQ),
.Q(CLBLL_L_X42Y68_SLICE_X68Y68_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLL_L_X42Y68_SLICE_X68Y68_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y80_SLICE_X69Y80_A5Q),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y68_SLICE_X68Y68_DO5),
.O6(CLBLL_L_X42Y68_SLICE_X68Y68_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f0f0f0f0)
  ) CLBLL_L_X42Y68_SLICE_X68Y68_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y80_SLICE_X69Y80_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y68_SLICE_X68Y68_CO5),
.O6(CLBLL_L_X42Y68_SLICE_X68Y68_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f0f0f0f0)
  ) CLBLL_L_X42Y68_SLICE_X68Y68_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y101_SLICE_X69Y101_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y68_SLICE_X68Y68_BO5),
.O6(CLBLL_L_X42Y68_SLICE_X68Y68_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff0000)
  ) CLBLL_L_X42Y68_SLICE_X68Y68_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X42Y80_SLICE_X69Y80_CQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y68_SLICE_X68Y68_AO5),
.O6(CLBLL_L_X42Y68_SLICE_X68Y68_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y68_SLICE_X69Y68_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y68_SLICE_X69Y68_DO5),
.O6(CLBLL_L_X42Y68_SLICE_X69Y68_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y68_SLICE_X69Y68_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y68_SLICE_X69Y68_CO5),
.O6(CLBLL_L_X42Y68_SLICE_X69Y68_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y68_SLICE_X69Y68_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y68_SLICE_X69Y68_BO5),
.O6(CLBLL_L_X42Y68_SLICE_X69Y68_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y68_SLICE_X69Y68_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y68_SLICE_X69Y68_AO5),
.O6(CLBLL_L_X42Y68_SLICE_X69Y68_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y69_SLICE_X68Y69_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y69_SLICE_X68Y69_AO5),
.Q(CLBLL_L_X42Y69_SLICE_X68Y69_AQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y69_SLICE_X68Y69_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y69_SLICE_X68Y69_BO5),
.Q(CLBLL_L_X42Y69_SLICE_X68Y69_BQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y69_SLICE_X68Y69_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y69_SLICE_X68Y69_CO5),
.Q(CLBLL_L_X42Y69_SLICE_X68Y69_CQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y69_SLICE_X68Y69_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y69_SLICE_X68Y69_DO5),
.Q(CLBLL_L_X42Y69_SLICE_X68Y69_DQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X42Y69_SLICE_X68Y69_CARRY4 (
.CI(1'b0),
.CO({CLBLL_L_X42Y69_SLICE_X68Y69_D_CY, CLBLL_L_X42Y69_SLICE_X68Y69_C_CY, CLBLL_L_X42Y69_SLICE_X68Y69_B_CY, CLBLL_L_X42Y69_SLICE_X68Y69_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({CLBLL_L_X42Y69_SLICE_X68Y69_D_XOR, CLBLL_L_X42Y69_SLICE_X68Y69_C_XOR, CLBLL_L_X42Y69_SLICE_X68Y69_B_XOR, CLBLL_L_X42Y69_SLICE_X68Y69_A_XOR}),
.S({CLBLL_L_X42Y69_SLICE_X68Y69_DO6, CLBLL_L_X42Y69_SLICE_X68Y69_CO6, CLBLL_L_X42Y69_SLICE_X68Y69_BO6, CLBLL_L_X42Y69_SLICE_X68Y69_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0f0f0f0)
  ) CLBLL_L_X42Y69_SLICE_X68Y69_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y70_SLICE_X68Y70_A_XOR),
.I3(1'b1),
.I4(CLBLL_L_X42Y70_SLICE_X68Y70_DQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y69_SLICE_X68Y69_DO5),
.O6(CLBLL_L_X42Y69_SLICE_X68Y69_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f0f0f0f0)
  ) CLBLL_L_X42Y69_SLICE_X68Y69_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y69_SLICE_X68Y69_B_XOR),
.I3(CLBLL_L_X42Y71_SLICE_X68Y71_B5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y69_SLICE_X68Y69_CO5),
.O6(CLBLL_L_X42Y69_SLICE_X68Y69_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLL_L_X42Y69_SLICE_X68Y69_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y69_SLICE_X68Y69_CQ),
.I2(1'b1),
.I3(CLBLL_L_X42Y70_SLICE_X68Y70_B_XOR),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y69_SLICE_X68Y69_BO5),
.O6(CLBLL_L_X42Y69_SLICE_X68Y69_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f00000ffff)
  ) CLBLL_L_X42Y69_SLICE_X68Y69_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y69_SLICE_X68Y69_AO5),
.I3(1'b1),
.I4(CLBLL_L_X42Y69_SLICE_X68Y69_AQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y69_SLICE_X68Y69_AO5),
.O6(CLBLL_L_X42Y69_SLICE_X68Y69_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y69_SLICE_X69Y69_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y69_SLICE_X69Y69_DO5),
.O6(CLBLL_L_X42Y69_SLICE_X69Y69_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000404)
  ) CLBLL_L_X42Y69_SLICE_X69Y69_CLUT (
.I0(CLBLL_L_X42Y69_SLICE_X68Y69_BQ),
.I1(CLBLL_L_X42Y71_SLICE_X68Y71_B5Q),
.I2(CLBLL_L_X42Y69_SLICE_X68Y69_DQ),
.I3(1'b1),
.I4(CLBLL_L_X42Y70_SLICE_X68Y70_DQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y69_SLICE_X69Y69_CO5),
.O6(CLBLL_L_X42Y69_SLICE_X69Y69_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y69_SLICE_X69Y69_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y69_SLICE_X69Y69_BO5),
.O6(CLBLL_L_X42Y69_SLICE_X69Y69_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y69_SLICE_X69Y69_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y69_SLICE_X69Y69_AO5),
.O6(CLBLL_L_X42Y69_SLICE_X69Y69_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y70_SLICE_X68Y70_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y70_SLICE_X68Y70_AO5),
.Q(CLBLL_L_X42Y70_SLICE_X68Y70_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y70_SLICE_X68Y70_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y71_SLICE_X68Y71_DO5),
.Q(CLBLL_L_X42Y70_SLICE_X68Y70_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y70_SLICE_X68Y70_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y70_SLICE_X68Y70_DO5),
.Q(CLBLL_L_X42Y70_SLICE_X68Y70_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X42Y70_SLICE_X68Y70_CARRY4 (
.CI(CLBLL_L_X42Y69_SLICE_X68Y69_COUT),
.CO({CLBLL_L_X42Y70_SLICE_X68Y70_COUT, CLBLL_L_X42Y70_SLICE_X68Y70_C_CY, CLBLL_L_X42Y70_SLICE_X68Y70_B_CY, CLBLL_L_X42Y70_SLICE_X68Y70_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, CLBLL_L_X42Y70_SLICE_X68Y70_BO5, 1'b0}),
.O({CLBLL_L_X42Y70_SLICE_X68Y70_D_XOR, CLBLL_L_X42Y70_SLICE_X68Y70_C_XOR, CLBLL_L_X42Y70_SLICE_X68Y70_B_XOR, CLBLL_L_X42Y70_SLICE_X68Y70_A_XOR}),
.S({CLBLL_L_X42Y70_SLICE_X68Y70_DO6, CLBLL_L_X42Y70_SLICE_X68Y70_CO6, CLBLL_L_X42Y70_SLICE_X68Y70_BO6, CLBLL_L_X42Y70_SLICE_X68Y70_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffff0000)
  ) CLBLL_L_X42Y70_SLICE_X68Y70_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y70_SLICE_X68Y70_BQ),
.I3(1'b1),
.I4(CLBLL_L_X42Y71_SLICE_X68Y71_BO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y70_SLICE_X68Y70_DO5),
.O6(CLBLL_L_X42Y70_SLICE_X68Y70_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLL_L_X42Y70_SLICE_X68Y70_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X42Y70_SLICE_X68Y70_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y70_SLICE_X68Y70_CO5),
.O6(CLBLL_L_X42Y70_SLICE_X68Y70_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaaaaaaa)
  ) CLBLL_L_X42Y70_SLICE_X68Y70_BLUT (
.I0(1'b0),
.I1(1'b1),
.I2(CLBLL_L_X42Y69_SLICE_X68Y69_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y70_SLICE_X68Y70_BO5),
.O6(CLBLL_L_X42Y70_SLICE_X68Y70_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaffff0000)
  ) CLBLL_L_X42Y70_SLICE_X68Y70_ALUT (
.I0(CLBLL_L_X42Y69_SLICE_X68Y69_DQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X42Y71_SLICE_X68Y71_DO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y70_SLICE_X68Y70_AO5),
.O6(CLBLL_L_X42Y70_SLICE_X68Y70_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y70_SLICE_X69Y70_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y70_SLICE_X69Y70_DO5),
.O6(CLBLL_L_X42Y70_SLICE_X69Y70_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y70_SLICE_X69Y70_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y70_SLICE_X69Y70_CO5),
.O6(CLBLL_L_X42Y70_SLICE_X69Y70_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y70_SLICE_X69Y70_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y70_SLICE_X69Y70_BO5),
.O6(CLBLL_L_X42Y70_SLICE_X69Y70_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y70_SLICE_X69Y70_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y70_SLICE_X69Y70_AO5),
.O6(CLBLL_L_X42Y70_SLICE_X69Y70_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y71_SLICE_X68Y71_B5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y69_SLICE_X68Y69_C_XOR),
.Q(CLBLL_L_X42Y71_SLICE_X68Y71_B5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y71_SLICE_X68Y71_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y71_SLICE_X68Y71_BO5),
.Q(CLBLL_L_X42Y71_SLICE_X68Y71_BQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h2200220022220000)
  ) CLBLL_L_X42Y71_SLICE_X68Y71_DLUT (
.I0(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I1(CLBLL_L_X42Y71_SLICE_X68Y71_CO5),
.I2(1'b1),
.I3(CLBLL_L_X42Y70_SLICE_X68Y70_C_XOR),
.I4(CLBLL_L_X42Y70_SLICE_X68Y70_D_XOR),
.I5(1'b1),
.O5(CLBLL_L_X42Y71_SLICE_X68Y71_DO5),
.O6(CLBLL_L_X42Y71_SLICE_X68Y71_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000022000000)
  ) CLBLL_L_X42Y71_SLICE_X68Y71_CLUT (
.I0(CLBLL_L_X42Y70_SLICE_X68Y70_AQ),
.I1(CLBLL_L_X42Y69_SLICE_X68Y69_C_XOR),
.I2(1'b1),
.I3(CLBLL_L_X42Y69_SLICE_X69Y69_CO5),
.I4(CLBLL_L_X42Y70_SLICE_X68Y70_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y71_SLICE_X68Y71_CO5),
.O6(CLBLL_L_X42Y71_SLICE_X68Y71_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h40404040aaaaaaaa)
  ) CLBLL_L_X42Y71_SLICE_X68Y71_BLUT (
.I0(CLBLL_L_X42Y71_SLICE_X68Y71_CO5),
.I1(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I2(CLBLL_L_X42Y69_SLICE_X68Y69_D_XOR),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y71_SLICE_X68Y71_BO5),
.O6(CLBLL_L_X42Y71_SLICE_X68Y71_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff887f0077007f00)
  ) CLBLL_L_X42Y71_SLICE_X68Y71_ALUT (
.I0(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I1(CLBLL_L_X42Y71_SLICE_X68Y71_BQ),
.I2(CLBLL_L_X42Y112_SLICE_X69Y112_DQ),
.I3(CLBLL_L_X42Y96_SLICE_X69Y96_B5Q),
.I4(CLBLL_L_X42Y112_SLICE_X69Y112_C5Q),
.I5(CLBLL_L_X42Y43_SLICE_X68Y43_B_XOR),
.O5(CLBLL_L_X42Y71_SLICE_X68Y71_AO5),
.O6(CLBLL_L_X42Y71_SLICE_X68Y71_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y71_SLICE_X69Y71_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y71_SLICE_X69Y71_DO5),
.O6(CLBLL_L_X42Y71_SLICE_X69Y71_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y71_SLICE_X69Y71_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y71_SLICE_X69Y71_CO5),
.O6(CLBLL_L_X42Y71_SLICE_X69Y71_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y71_SLICE_X69Y71_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y71_SLICE_X69Y71_BO5),
.O6(CLBLL_L_X42Y71_SLICE_X69Y71_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y71_SLICE_X69Y71_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y71_SLICE_X69Y71_AO5),
.O6(CLBLL_L_X42Y71_SLICE_X69Y71_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y80_SLICE_X68Y80_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y80_SLICE_X68Y80_DO5),
.O6(CLBLL_L_X42Y80_SLICE_X68Y80_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y80_SLICE_X68Y80_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y80_SLICE_X68Y80_CO5),
.O6(CLBLL_L_X42Y80_SLICE_X68Y80_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y80_SLICE_X68Y80_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y80_SLICE_X68Y80_BO5),
.O6(CLBLL_L_X42Y80_SLICE_X68Y80_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y80_SLICE_X68Y80_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y80_SLICE_X68Y80_AO5),
.O6(CLBLL_L_X42Y80_SLICE_X68Y80_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y80_SLICE_X69Y80_A5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y96_SLICE_X68Y96_DQ),
.Q(CLBLL_L_X42Y80_SLICE_X69Y80_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y80_SLICE_X69Y80_B5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(BRAM_L_X44Y95_RAMB18_X2Y38_DO0),
.Q(CLBLL_L_X42Y80_SLICE_X69Y80_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y80_SLICE_X69Y80_C5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y92_SLICE_X69Y92_DQ),
.Q(CLBLL_L_X42Y80_SLICE_X69Y80_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y80_SLICE_X69Y80_D5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y93_SLICE_X68Y93_A5Q),
.Q(CLBLL_L_X42Y80_SLICE_X69Y80_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y80_SLICE_X69Y80_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y80_SLICE_X69Y80_AO5),
.Q(CLBLL_L_X42Y80_SLICE_X69Y80_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y80_SLICE_X69Y80_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y80_SLICE_X69Y80_BO5),
.Q(CLBLL_L_X42Y80_SLICE_X69Y80_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y80_SLICE_X69Y80_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y80_SLICE_X69Y80_CO5),
.Q(CLBLL_L_X42Y80_SLICE_X69Y80_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y80_SLICE_X69Y80_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y80_SLICE_X69Y80_DO5),
.Q(CLBLL_L_X42Y80_SLICE_X69Y80_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLL_L_X42Y80_SLICE_X69Y80_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y96_SLICE_X68Y96_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y80_SLICE_X69Y80_DO5),
.O6(CLBLL_L_X42Y80_SLICE_X69Y80_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLL_L_X42Y80_SLICE_X69Y80_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_L_X44Y95_RAMB18_X2Y38_DO13),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y80_SLICE_X69Y80_CO5),
.O6(CLBLL_L_X42Y80_SLICE_X69Y80_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff0000)
  ) CLBLL_L_X42Y80_SLICE_X69Y80_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(BRAM_L_X44Y95_RAMB18_X2Y38_DO1),
.I5(1'b1),
.O5(CLBLL_L_X42Y80_SLICE_X69Y80_BO5),
.O6(CLBLL_L_X42Y80_SLICE_X69Y80_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLL_L_X42Y80_SLICE_X69Y80_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_L_X44Y95_RAMB18_X2Y38_DO3),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y80_SLICE_X69Y80_AO5),
.O6(CLBLL_L_X42Y80_SLICE_X69Y80_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y90_SLICE_X68Y90_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y90_SLICE_X68Y90_AO5),
.Q(CLBLL_L_X42Y90_SLICE_X68Y90_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y90_SLICE_X68Y90_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y90_SLICE_X68Y90_BO5),
.Q(CLBLL_L_X42Y90_SLICE_X68Y90_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y90_SLICE_X68Y90_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y90_SLICE_X68Y90_DO5),
.Q(CLBLL_L_X42Y90_SLICE_X68Y90_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X42Y90_SLICE_X68Y90_CARRY4 (
.CI(1'b0),
.CO({CLBLL_L_X42Y90_SLICE_X68Y90_D_CY, CLBLL_L_X42Y90_SLICE_X68Y90_C_CY, CLBLL_L_X42Y90_SLICE_X68Y90_B_CY, CLBLL_L_X42Y90_SLICE_X68Y90_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({CLBLL_L_X42Y90_SLICE_X68Y90_D_XOR, CLBLL_L_X42Y90_SLICE_X68Y90_C_XOR, CLBLL_L_X42Y90_SLICE_X68Y90_B_XOR, CLBLL_L_X42Y90_SLICE_X68Y90_A_XOR}),
.S({CLBLL_L_X42Y90_SLICE_X68Y90_DO6, CLBLL_L_X42Y90_SLICE_X68Y90_CO6, CLBLL_L_X42Y90_SLICE_X68Y90_BO6, CLBLL_L_X42Y90_SLICE_X68Y90_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_L_X42Y90_SLICE_X68Y90_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y90_SLICE_X69Y90_DO6),
.I2(CLBLL_L_X42Y90_SLICE_X68Y90_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y90_SLICE_X68Y90_DO5),
.O6(CLBLL_L_X42Y90_SLICE_X68Y90_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLL_L_X42Y90_SLICE_X68Y90_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y90_SLICE_X68Y90_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y90_SLICE_X68Y90_CO5),
.O6(CLBLL_L_X42Y90_SLICE_X68Y90_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLL_L_X42Y90_SLICE_X68Y90_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y90_SLICE_X68Y90_BQ),
.I2(1'b1),
.I3(CLBLL_L_X42Y90_SLICE_X69Y90_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y90_SLICE_X68Y90_BO5),
.O6(CLBLL_L_X42Y90_SLICE_X68Y90_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_L_X42Y90_SLICE_X68Y90_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y90_SLICE_X69Y90_BO5),
.I2(CLBLL_L_X42Y91_SLICE_X69Y91_AO5),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y90_SLICE_X68Y90_AO5),
.O6(CLBLL_L_X42Y90_SLICE_X68Y90_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y90_SLICE_X69Y90_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y96_SLICE_X68Y96_AO6),
.D(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.Q(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf777800000000000)
  ) CLBLL_L_X42Y90_SLICE_X69Y90_DLUT (
.I0(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I1(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I2(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I3(CLBLL_L_X42Y90_SLICE_X68Y90_C_XOR),
.I4(CLBLL_L_X42Y90_SLICE_X68Y90_DQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y90_SLICE_X69Y90_DO5),
.O6(CLBLL_L_X42Y90_SLICE_X69Y90_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf870707000000000)
  ) CLBLL_L_X42Y90_SLICE_X69Y90_CLUT (
.I0(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I1(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I2(CLBLL_L_X42Y90_SLICE_X68Y90_BQ),
.I3(CLBLL_L_X42Y90_SLICE_X68Y90_B_XOR),
.I4(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y90_SLICE_X69Y90_CO5),
.O6(CLBLL_L_X42Y90_SLICE_X69Y90_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000088f0f0f0)
  ) CLBLL_L_X42Y90_SLICE_X69Y90_BLUT (
.I0(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I1(CLBLL_L_X42Y90_SLICE_X68Y90_D_XOR),
.I2(CLBLL_L_X42Y90_SLICE_X68Y90_AQ),
.I3(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I4(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y90_SLICE_X69Y90_BO5),
.O6(CLBLL_L_X42Y90_SLICE_X69Y90_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000e2aa22aa)
  ) CLBLL_L_X42Y90_SLICE_X69Y90_ALUT (
.I0(CLBLL_L_X42Y91_SLICE_X68Y91_AQ),
.I1(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I2(CLBLL_L_X42Y91_SLICE_X68Y91_A_XOR),
.I3(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I4(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y90_SLICE_X69Y90_AO5),
.O6(CLBLL_L_X42Y90_SLICE_X69Y90_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y91_SLICE_X68Y91_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y91_SLICE_X68Y91_AO5),
.Q(CLBLL_L_X42Y91_SLICE_X68Y91_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y91_SLICE_X68Y91_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y91_SLICE_X68Y91_BO5),
.Q(CLBLL_L_X42Y91_SLICE_X68Y91_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y91_SLICE_X68Y91_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y91_SLICE_X68Y91_CO5),
.Q(CLBLL_L_X42Y91_SLICE_X68Y91_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y91_SLICE_X68Y91_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y91_SLICE_X68Y91_DO5),
.Q(CLBLL_L_X42Y91_SLICE_X68Y91_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X42Y91_SLICE_X68Y91_CARRY4 (
.CI(CLBLL_L_X42Y90_SLICE_X68Y90_COUT),
.CO({CLBLL_L_X42Y91_SLICE_X68Y91_COUT, CLBLL_L_X42Y91_SLICE_X68Y91_C_CY, CLBLL_L_X42Y91_SLICE_X68Y91_B_CY, CLBLL_L_X42Y91_SLICE_X68Y91_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_L_X42Y91_SLICE_X68Y91_D_XOR, CLBLL_L_X42Y91_SLICE_X68Y91_C_XOR, CLBLL_L_X42Y91_SLICE_X68Y91_B_XOR, CLBLL_L_X42Y91_SLICE_X68Y91_A_XOR}),
.S({CLBLL_L_X42Y91_SLICE_X68Y91_DO6, CLBLL_L_X42Y91_SLICE_X68Y91_CO6, CLBLL_L_X42Y91_SLICE_X68Y91_BO6, CLBLL_L_X42Y91_SLICE_X68Y91_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ff00)
  ) CLBLL_L_X42Y91_SLICE_X68Y91_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y91_SLICE_X68Y91_DQ),
.I3(CLBLL_L_X42Y94_SLICE_X69Y94_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y91_SLICE_X68Y91_DO5),
.O6(CLBLL_L_X42Y91_SLICE_X68Y91_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLL_L_X42Y91_SLICE_X68Y91_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y91_SLICE_X68Y91_CQ),
.I2(1'b1),
.I3(CLBLL_L_X42Y94_SLICE_X69Y94_BO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y91_SLICE_X68Y91_CO5),
.O6(CLBLL_L_X42Y91_SLICE_X68Y91_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLL_L_X42Y91_SLICE_X68Y91_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y91_SLICE_X68Y91_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X42Y94_SLICE_X69Y94_DO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y91_SLICE_X68Y91_BO5),
.O6(CLBLL_L_X42Y91_SLICE_X68Y91_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLL_L_X42Y91_SLICE_X68Y91_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y91_SLICE_X68Y91_AQ),
.I2(1'b1),
.I3(CLBLL_L_X42Y90_SLICE_X69Y90_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y91_SLICE_X68Y91_AO5),
.O6(CLBLL_L_X42Y91_SLICE_X68Y91_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y91_SLICE_X69Y91_D5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y91_SLICE_X69Y91_DQ),
.Q(CLBLL_L_X42Y91_SLICE_X69Y91_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y91_SLICE_X69Y91_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y91_SLICE_X69Y91_BQ),
.Q(CLBLL_L_X42Y91_SLICE_X69Y91_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y91_SLICE_X69Y91_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y91_SLICE_X69Y91_BO5),
.Q(CLBLL_L_X42Y91_SLICE_X69Y91_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y91_SLICE_X69Y91_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y91_SLICE_X69Y91_CO6),
.Q(CLBLL_L_X42Y91_SLICE_X69Y91_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y91_SLICE_X69Y91_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y91_SLICE_X69Y91_DO5),
.Q(CLBLL_L_X42Y91_SLICE_X69Y91_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000c0aaaaaa)
  ) CLBLL_L_X42Y91_SLICE_X69Y91_DLUT (
.I0(CLBLL_L_X42Y91_SLICE_X69Y91_DQ),
.I1(CLBLL_L_X42Y94_SLICE_X68Y94_B_XOR),
.I2(CLBLL_L_X42Y96_SLICE_X68Y96_AO5),
.I3(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I4(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y91_SLICE_X69Y91_DO5),
.O6(CLBLL_L_X42Y91_SLICE_X69Y91_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf5f800000000000)
  ) CLBLL_L_X42Y91_SLICE_X69Y91_CLUT (
.I0(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I1(CLBLL_L_X42Y96_SLICE_X68Y96_AO5),
.I2(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I3(CLBLL_L_X42Y94_SLICE_X68Y94_C_XOR),
.I4(CLBLL_L_X42Y91_SLICE_X69Y91_CQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y91_SLICE_X69Y91_CO5),
.O6(CLBLL_L_X42Y91_SLICE_X69Y91_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000e222aaaa)
  ) CLBLL_L_X42Y91_SLICE_X69Y91_BLUT (
.I0(CLBLL_L_X42Y91_SLICE_X69Y91_BQ),
.I1(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I2(CLBLL_L_X42Y96_SLICE_X68Y96_AO5),
.I3(CLBLL_L_X42Y93_SLICE_X68Y93_D_XOR),
.I4(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y91_SLICE_X69Y91_BO5),
.O6(CLBLL_L_X42Y91_SLICE_X69Y91_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h777788000000ffff)
  ) CLBLL_L_X42Y91_SLICE_X69Y91_ALUT (
.I0(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I1(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I2(1'b1),
.I3(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I4(CLBLL_L_X42Y94_SLICE_X68Y94_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y91_SLICE_X69Y91_AO5),
.O6(CLBLL_L_X42Y91_SLICE_X69Y91_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y92_SLICE_X68Y92_D5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y92_SLICE_X69Y92_C5Q),
.Q(CLBLL_L_X42Y92_SLICE_X68Y92_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y92_SLICE_X68Y92_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y92_SLICE_X68Y92_AO5),
.Q(CLBLL_L_X42Y92_SLICE_X68Y92_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y92_SLICE_X68Y92_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y92_SLICE_X68Y92_BO5),
.Q(CLBLL_L_X42Y92_SLICE_X68Y92_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y92_SLICE_X68Y92_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y92_SLICE_X68Y92_CO5),
.Q(CLBLL_L_X42Y92_SLICE_X68Y92_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X42Y92_SLICE_X68Y92_CARRY4 (
.CI(CLBLL_L_X42Y91_SLICE_X68Y91_COUT),
.CO({CLBLL_L_X42Y92_SLICE_X68Y92_COUT, CLBLL_L_X42Y92_SLICE_X68Y92_C_CY, CLBLL_L_X42Y92_SLICE_X68Y92_B_CY, CLBLL_L_X42Y92_SLICE_X68Y92_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_L_X42Y92_SLICE_X68Y92_DO5, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_L_X42Y92_SLICE_X68Y92_D_XOR, CLBLL_L_X42Y92_SLICE_X68Y92_C_XOR, CLBLL_L_X42Y92_SLICE_X68Y92_B_XOR, CLBLL_L_X42Y92_SLICE_X68Y92_A_XOR}),
.S({CLBLL_L_X42Y92_SLICE_X68Y92_DO6, CLBLL_L_X42Y92_SLICE_X68Y92_CO6, CLBLL_L_X42Y92_SLICE_X68Y92_BO6, CLBLL_L_X42Y92_SLICE_X68Y92_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccccccccccc)
  ) CLBLL_L_X42Y92_SLICE_X68Y92_DLUT (
.I0(1'b1),
.I1(1'b0),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y92_SLICE_X68Y92_DO5),
.O6(CLBLL_L_X42Y92_SLICE_X68Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ff00)
  ) CLBLL_L_X42Y92_SLICE_X68Y92_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b0),
.I3(BRAM_L_X44Y95_RAMB18_X2Y38_DO14),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y92_SLICE_X68Y92_CO5),
.O6(CLBLL_L_X42Y92_SLICE_X68Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLL_L_X42Y92_SLICE_X68Y92_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y92_SLICE_X69Y92_AQ),
.I2(CLBLL_L_X42Y92_SLICE_X69Y92_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y92_SLICE_X68Y92_BO5),
.O6(CLBLL_L_X42Y92_SLICE_X68Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00cccccccc)
  ) CLBLL_L_X42Y92_SLICE_X68Y92_ALUT (
.I0(1'b1),
.I1(BRAM_L_X44Y95_RAMB18_X2Y38_DO12),
.I2(1'b1),
.I3(CLBLL_L_X42Y92_SLICE_X69Y92_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y92_SLICE_X68Y92_AO5),
.O6(CLBLL_L_X42Y92_SLICE_X68Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y92_SLICE_X69Y92_B5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y92_SLICE_X69Y92_BO5),
.Q(CLBLL_L_X42Y92_SLICE_X69Y92_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y92_SLICE_X69Y92_C5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y92_SLICE_X69Y92_CO5),
.Q(CLBLL_L_X42Y92_SLICE_X69Y92_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y92_SLICE_X69Y92_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y92_SLICE_X69Y92_AO5),
.Q(CLBLL_L_X42Y92_SLICE_X69Y92_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y92_SLICE_X69Y92_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y92_SLICE_X69Y92_AO6),
.Q(CLBLL_L_X42Y92_SLICE_X69Y92_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y92_SLICE_X69Y92_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y92_SLICE_X69Y92_DO5),
.Q(CLBLL_L_X42Y92_SLICE_X69Y92_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000008f80ff00)
  ) CLBLL_L_X42Y92_SLICE_X69Y92_DLUT (
.I0(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I1(CLBLL_L_X42Y92_SLICE_X68Y92_B_XOR),
.I2(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I3(CLBLL_L_X42Y92_SLICE_X69Y92_DQ),
.I4(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y92_SLICE_X69Y92_DO5),
.O6(CLBLL_L_X42Y92_SLICE_X69Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000c0aaaaaa)
  ) CLBLL_L_X42Y92_SLICE_X69Y92_CLUT (
.I0(CLBLL_L_X42Y92_SLICE_X69Y92_C5Q),
.I1(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I2(CLBLL_L_X42Y92_SLICE_X68Y92_A_XOR),
.I3(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I4(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y92_SLICE_X69Y92_CO5),
.O6(CLBLL_L_X42Y92_SLICE_X69Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000005fa0ff00)
  ) CLBLL_L_X42Y92_SLICE_X69Y92_BLUT (
.I0(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I1(1'b1),
.I2(CLBLL_L_X42Y95_SLICE_X68Y95_D5Q),
.I3(CLBLL_L_X42Y92_SLICE_X69Y92_B5Q),
.I4(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y92_SLICE_X69Y92_BO5),
.O6(CLBLL_L_X42Y92_SLICE_X69Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hd5ff8000ffff0000)
  ) CLBLL_L_X42Y92_SLICE_X69Y92_ALUT (
.I0(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I1(CLBLL_L_X42Y94_SLICE_X68Y94_A_XOR),
.I2(CLBLL_L_X42Y96_SLICE_X68Y96_AO5),
.I3(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I4(CLBLL_L_X42Y92_SLICE_X69Y92_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y92_SLICE_X69Y92_AO5),
.O6(CLBLL_L_X42Y92_SLICE_X69Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y93_SLICE_X68Y93_A5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.D(CLBLL_L_X42Y93_SLICE_X68Y93_AO5),
.Q(CLBLL_L_X42Y93_SLICE_X68Y93_A5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y93_SLICE_X68Y93_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.D(1'b0),
.Q(CLBLL_L_X42Y93_SLICE_X68Y93_BQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y93_SLICE_X68Y93_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.D(1'b0),
.Q(CLBLL_L_X42Y93_SLICE_X68Y93_CQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y93_SLICE_X68Y93_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.D(1'b0),
.Q(CLBLL_L_X42Y93_SLICE_X68Y93_DQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X42Y93_SLICE_X68Y93_CARRY4 (
.CI(1'b0),
.CO({CLBLL_L_X42Y93_SLICE_X68Y93_D_CY, CLBLL_L_X42Y93_SLICE_X68Y93_C_CY, CLBLL_L_X42Y93_SLICE_X68Y93_B_CY, CLBLL_L_X42Y93_SLICE_X68Y93_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({CLBLL_L_X42Y93_SLICE_X68Y93_D_XOR, CLBLL_L_X42Y93_SLICE_X68Y93_C_XOR, CLBLL_L_X42Y93_SLICE_X68Y93_B_XOR, CLBLL_L_X42Y93_SLICE_X68Y93_A_XOR}),
.S({CLBLL_L_X42Y93_SLICE_X68Y93_DO6, CLBLL_L_X42Y93_SLICE_X68Y93_CO6, CLBLL_L_X42Y93_SLICE_X68Y93_BO6, CLBLL_L_X42Y93_SLICE_X68Y93_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000000000)
  ) CLBLL_L_X42Y93_SLICE_X68Y93_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X42Y91_SLICE_X69Y91_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y93_SLICE_X68Y93_DO5),
.O6(CLBLL_L_X42Y93_SLICE_X68Y93_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLL_L_X42Y93_SLICE_X68Y93_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X42Y95_SLICE_X69Y95_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y93_SLICE_X68Y93_CO5),
.O6(CLBLL_L_X42Y93_SLICE_X68Y93_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLL_L_X42Y93_SLICE_X68Y93_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y97_SLICE_X68Y97_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y93_SLICE_X68Y93_BO5),
.O6(CLBLL_L_X42Y93_SLICE_X68Y93_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f05555ffff)
  ) CLBLL_L_X42Y93_SLICE_X68Y93_ALUT (
.I0(CLBLL_L_X42Y92_SLICE_X68Y92_C_XOR),
.I1(1'b1),
.I2(CLBLL_L_X42Y96_SLICE_X68Y96_BO5),
.I3(1'b1),
.I4(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y93_SLICE_X68Y93_AO5),
.O6(CLBLL_L_X42Y93_SLICE_X68Y93_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y93_SLICE_X69Y93_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y91_SLICE_X69Y91_CQ),
.Q(CLBLL_L_X42Y93_SLICE_X69Y93_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf500310000000000)
  ) CLBLL_L_X42Y93_SLICE_X69Y93_DLUT (
.I0(CLBLL_L_X42Y92_SLICE_X69Y92_AQ),
.I1(CLBLL_L_X42Y96_SLICE_X68Y96_AQ),
.I2(BRAM_L_X44Y95_RAMB18_X2Y38_DO4),
.I3(CLBLL_L_X42Y93_SLICE_X69Y93_BO5),
.I4(BRAM_L_X44Y95_RAMB18_X2Y38_DO0),
.I5(1'b1),
.O5(CLBLL_L_X42Y93_SLICE_X69Y93_DO5),
.O6(CLBLL_L_X42Y93_SLICE_X69Y93_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000084000000)
  ) CLBLL_L_X42Y93_SLICE_X69Y93_CLUT (
.I0(CLBLL_L_X42Y96_SLICE_X68Y96_DQ),
.I1(CLBLL_L_X42Y93_SLICE_X69Y93_AO6),
.I2(BRAM_L_X44Y95_RAMB18_X2Y38_DO8),
.I3(CLBLL_L_X42Y93_SLICE_X69Y93_DO6),
.I4(CLBLL_L_X42Y95_SLICE_X68Y95_CO5),
.I5(1'b1),
.O5(CLBLL_L_X42Y93_SLICE_X69Y93_CO5),
.O6(CLBLL_L_X42Y93_SLICE_X69Y93_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000003)
  ) CLBLL_L_X42Y93_SLICE_X69Y93_BLUT (
.I0(1'b1),
.I1(BRAM_L_X44Y95_RAMB18_X2Y38_DO11),
.I2(BRAM_L_X44Y95_RAMB18_X2Y38_DO14),
.I3(BRAM_L_X44Y95_RAMB18_X2Y38_DO13),
.I4(BRAM_L_X44Y95_RAMB18_X2Y38_DO12),
.I5(1'b1),
.O5(CLBLL_L_X42Y93_SLICE_X69Y93_BO5),
.O6(CLBLL_L_X42Y93_SLICE_X69Y93_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h8200410000820041)
  ) CLBLL_L_X42Y93_SLICE_X69Y93_ALUT (
.I0(CLBLL_L_X42Y91_SLICE_X69Y91_AQ),
.I1(CLBLL_L_X42Y93_SLICE_X69Y93_BQ),
.I2(BRAM_L_X44Y95_RAMB18_X2Y38_DO6),
.I3(BRAM_L_X44Y95_RAMB18_X2Y38_DO1),
.I4(BRAM_L_X44Y95_RAMB18_X2Y38_DO3),
.I5(CLBLL_L_X42Y97_SLICE_X68Y97_AQ),
.O5(CLBLL_L_X42Y93_SLICE_X69Y93_AO5),
.O6(CLBLL_L_X42Y93_SLICE_X69Y93_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y94_SLICE_X68Y94_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y94_SLICE_X68Y94_BO5),
.Q(CLBLL_L_X42Y94_SLICE_X68Y94_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X42Y94_SLICE_X68Y94_CARRY4 (
.CI(CLBLL_L_X42Y93_SLICE_X68Y93_COUT),
.CO({CLBLL_L_X42Y94_SLICE_X68Y94_COUT, CLBLL_L_X42Y94_SLICE_X68Y94_C_CY, CLBLL_L_X42Y94_SLICE_X68Y94_B_CY, CLBLL_L_X42Y94_SLICE_X68Y94_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_L_X42Y94_SLICE_X68Y94_D_XOR, CLBLL_L_X42Y94_SLICE_X68Y94_C_XOR, CLBLL_L_X42Y94_SLICE_X68Y94_B_XOR, CLBLL_L_X42Y94_SLICE_X68Y94_A_XOR}),
.S({CLBLL_L_X42Y94_SLICE_X68Y94_DO6, CLBLL_L_X42Y94_SLICE_X68Y94_CO6, CLBLL_L_X42Y94_SLICE_X68Y94_BO6, CLBLL_L_X42Y94_SLICE_X68Y94_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000000000)
  ) CLBLL_L_X42Y94_SLICE_X68Y94_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X42Y95_SLICE_X69Y95_DQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y94_SLICE_X68Y94_DO5),
.O6(CLBLL_L_X42Y94_SLICE_X68Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLL_L_X42Y94_SLICE_X68Y94_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X42Y91_SLICE_X69Y91_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y94_SLICE_X68Y94_CO5),
.O6(CLBLL_L_X42Y94_SLICE_X68Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaaaaaaa)
  ) CLBLL_L_X42Y94_SLICE_X68Y94_BLUT (
.I0(CLBLL_L_X42Y91_SLICE_X69Y91_AO6),
.I1(1'b1),
.I2(CLBLL_L_X42Y91_SLICE_X69Y91_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y94_SLICE_X68Y94_BO5),
.O6(CLBLL_L_X42Y94_SLICE_X68Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLL_L_X42Y94_SLICE_X68Y94_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y92_SLICE_X69Y92_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y94_SLICE_X68Y94_AO5),
.O6(CLBLL_L_X42Y94_SLICE_X68Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y94_SLICE_X69Y94_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(1'b1),
.Q(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'he222aaaa00000000)
  ) CLBLL_L_X42Y94_SLICE_X69Y94_DLUT (
.I0(CLBLL_L_X42Y91_SLICE_X68Y91_BQ),
.I1(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I2(CLBLL_L_X42Y91_SLICE_X68Y91_B_XOR),
.I3(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I4(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y94_SLICE_X69Y94_DO5),
.O6(CLBLL_L_X42Y94_SLICE_X69Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y94_SLICE_X69Y94_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y94_SLICE_X69Y94_CO5),
.O6(CLBLL_L_X42Y94_SLICE_X69Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000e2aa22aa)
  ) CLBLL_L_X42Y94_SLICE_X69Y94_BLUT (
.I0(CLBLL_L_X42Y91_SLICE_X68Y91_CQ),
.I1(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I2(CLBLL_L_X42Y91_SLICE_X68Y91_C_XOR),
.I3(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I4(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y94_SLICE_X69Y94_BO5),
.O6(CLBLL_L_X42Y94_SLICE_X69Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000008f80ff00)
  ) CLBLL_L_X42Y94_SLICE_X69Y94_ALUT (
.I0(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I1(CLBLL_L_X42Y91_SLICE_X68Y91_D_XOR),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(CLBLL_L_X42Y91_SLICE_X68Y91_DQ),
.I4(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y94_SLICE_X69Y94_AO5),
.O6(CLBLL_L_X42Y94_SLICE_X69Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y95_SLICE_X68Y95_D5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y95_SLICE_X69Y95_AO6),
.Q(CLBLL_L_X42Y95_SLICE_X68Y95_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X42Y95_SLICE_X68Y95_CARRY4 (
.CI(CLBLL_L_X42Y94_SLICE_X68Y94_COUT),
.CO({CLBLL_L_X42Y95_SLICE_X68Y95_COUT, CLBLL_L_X42Y95_SLICE_X68Y95_C_CY, CLBLL_L_X42Y95_SLICE_X68Y95_B_CY, CLBLL_L_X42Y95_SLICE_X68Y95_A_CY}),
.CYINIT(1'b0),
.DI({CLBLL_L_X42Y95_SLICE_X68Y95_DO5, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_L_X42Y95_SLICE_X68Y95_D_XOR, CLBLL_L_X42Y95_SLICE_X68Y95_C_XOR, CLBLL_L_X42Y95_SLICE_X68Y95_B_XOR, CLBLL_L_X42Y95_SLICE_X68Y95_A_XOR}),
.S({CLBLL_L_X42Y95_SLICE_X68Y95_DO6, CLBLL_L_X42Y95_SLICE_X68Y95_CO6, CLBLL_L_X42Y95_SLICE_X68Y95_BO6, CLBLL_L_X42Y95_SLICE_X68Y95_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccccccccccc)
  ) CLBLL_L_X42Y95_SLICE_X68Y95_DLUT (
.I0(1'b1),
.I1(1'b0),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y95_SLICE_X68Y95_DO5),
.O6(CLBLL_L_X42Y95_SLICE_X68Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0bbbb00bb)
  ) CLBLL_L_X42Y95_SLICE_X68Y95_CLUT (
.I0(CLBLL_L_X42Y96_SLICE_X68Y96_AQ),
.I1(BRAM_L_X44Y95_RAMB18_X2Y38_DO0),
.I2(1'b0),
.I3(CLBLL_L_X42Y95_SLICE_X69Y95_D5Q),
.I4(BRAM_L_X44Y95_RAMB18_X2Y38_DO7),
.I5(1'b1),
.O5(CLBLL_L_X42Y95_SLICE_X68Y95_CO5),
.O6(CLBLL_L_X42Y95_SLICE_X68Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLL_L_X42Y95_SLICE_X68Y95_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y96_SLICE_X68Y96_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y95_SLICE_X68Y95_BO5),
.O6(CLBLL_L_X42Y95_SLICE_X68Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000000000)
  ) CLBLL_L_X42Y95_SLICE_X68Y95_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X42Y95_SLICE_X69Y95_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X42Y95_SLICE_X68Y95_AO5),
.O6(CLBLL_L_X42Y95_SLICE_X68Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y95_SLICE_X69Y95_A5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y95_SLICE_X69Y95_CO6),
.Q(CLBLL_L_X42Y95_SLICE_X69Y95_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y95_SLICE_X69Y95_D5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y95_SLICE_X69Y95_DQ),
.Q(CLBLL_L_X42Y95_SLICE_X69Y95_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y95_SLICE_X69Y95_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y95_SLICE_X69Y95_AO5),
.Q(CLBLL_L_X42Y95_SLICE_X69Y95_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y95_SLICE_X69Y95_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y95_SLICE_X69Y95_BO5),
.Q(CLBLL_L_X42Y95_SLICE_X69Y95_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y95_SLICE_X69Y95_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y95_SLICE_X69Y95_CO5),
.Q(CLBLL_L_X42Y95_SLICE_X69Y95_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y95_SLICE_X69Y95_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y95_SLICE_X69Y95_DO5),
.Q(CLBLL_L_X42Y95_SLICE_X69Y95_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f7807700)
  ) CLBLL_L_X42Y95_SLICE_X69Y95_DLUT (
.I0(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I1(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I2(CLBLL_L_X42Y96_SLICE_X68Y96_AO5),
.I3(CLBLL_L_X42Y95_SLICE_X69Y95_DQ),
.I4(CLBLL_L_X42Y94_SLICE_X68Y94_D_XOR),
.I5(1'b1),
.O5(CLBLL_L_X42Y95_SLICE_X69Y95_DO5),
.O6(CLBLL_L_X42Y95_SLICE_X69Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7807700ff00ff00)
  ) CLBLL_L_X42Y95_SLICE_X69Y95_CLUT (
.I0(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I1(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I2(CLBLL_L_X42Y96_SLICE_X68Y96_AO5),
.I3(CLBLL_L_X42Y95_SLICE_X69Y95_A5Q),
.I4(CLBLL_L_X42Y95_SLICE_X68Y95_A_XOR),
.I5(1'b1),
.O5(CLBLL_L_X42Y95_SLICE_X69Y95_CO5),
.O6(CLBLL_L_X42Y95_SLICE_X69Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f7807700)
  ) CLBLL_L_X42Y95_SLICE_X69Y95_BLUT (
.I0(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I1(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I2(CLBLL_L_X42Y93_SLICE_X68Y93_C_XOR),
.I3(CLBLL_L_X42Y95_SLICE_X69Y95_BQ),
.I4(CLBLL_L_X42Y96_SLICE_X68Y96_AO5),
.I5(1'b1),
.O5(CLBLL_L_X42Y95_SLICE_X69Y95_BO5),
.O6(CLBLL_L_X42Y95_SLICE_X69Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5af05af0ffff0000)
  ) CLBLL_L_X42Y95_SLICE_X69Y95_ALUT (
.I0(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I1(1'b1),
.I2(CLBLL_L_X42Y95_SLICE_X68Y95_D5Q),
.I3(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I4(CLBLL_L_X42Y95_SLICE_X69Y95_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y95_SLICE_X69Y95_AO5),
.O6(CLBLL_L_X42Y95_SLICE_X69Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y96_SLICE_X68Y96_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y96_SLICE_X68Y96_BQ),
.Q(CLBLL_L_X42Y96_SLICE_X68Y96_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y96_SLICE_X68Y96_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y96_SLICE_X68Y96_CO6),
.Q(CLBLL_L_X42Y96_SLICE_X68Y96_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y96_SLICE_X68Y96_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y96_SLICE_X68Y96_DO5),
.Q(CLBLL_L_X42Y96_SLICE_X68Y96_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y96_SLICE_X68Y96_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y96_SLICE_X68Y96_CQ),
.Q(CLBLL_L_X42Y96_SLICE_X68Y96_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000caaa0aaa)
  ) CLBLL_L_X42Y96_SLICE_X68Y96_DLUT (
.I0(CLBLL_L_X42Y96_SLICE_X68Y96_CQ),
.I1(CLBLL_L_X42Y95_SLICE_X68Y95_B_XOR),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I4(CLBLL_L_X42Y96_SLICE_X68Y96_AO5),
.I5(1'b1),
.O5(CLBLL_L_X42Y96_SLICE_X68Y96_DO5),
.O6(CLBLL_L_X42Y96_SLICE_X68Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h777780800a0a0a0a)
  ) CLBLL_L_X42Y96_SLICE_X68Y96_CLUT (
.I0(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I1(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I2(CLBLL_L_X42Y96_SLICE_X68Y96_AO5),
.I3(1'b1),
.I4(CLBLL_L_X42Y96_SLICE_X68Y96_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y96_SLICE_X68Y96_CO5),
.O6(CLBLL_L_X42Y96_SLICE_X68Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h222200000f0f0f0f)
  ) CLBLL_L_X42Y96_SLICE_X68Y96_BLUT (
.I0(CLBLL_L_X42Y97_SLICE_X68Y97_DO5),
.I1(CLBLL_L_X42Y113_SLICE_X68Y113_D5Q),
.I2(CLBLL_L_X42Y96_SLICE_X68Y96_BQ),
.I3(1'b1),
.I4(CLBLL_L_X42Y93_SLICE_X68Y93_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X42Y96_SLICE_X68Y96_BO5),
.O6(CLBLL_L_X42Y96_SLICE_X68Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555000000f000f0)
  ) CLBLL_L_X42Y96_SLICE_X68Y96_ALUT (
.I0(CLBLL_L_X42Y96_SLICE_X68Y96_AO5),
.I1(1'b1),
.I2(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I3(CLBLL_L_X42Y92_SLICE_X68Y92_C_XOR),
.I4(CLBLL_L_X42Y96_SLICE_X68Y96_DO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y96_SLICE_X68Y96_AO5),
.O6(CLBLL_L_X42Y96_SLICE_X68Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y96_SLICE_X69Y96_B5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y71_SLICE_X68Y71_AO6),
.Q(CLBLL_L_X42Y96_SLICE_X69Y96_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y96_SLICE_X69Y96_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y96_SLICE_X69Y96_BO5),
.Q(CLBLL_L_X42Y96_SLICE_X69Y96_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hdf8fd585da8ad080)
  ) CLBLL_L_X42Y96_SLICE_X69Y96_DLUT (
.I0(CLBLL_L_X42Y96_SLICE_X69Y96_BQ),
.I1(CLBLL_L_X42Y118_SLICE_X69Y118_DQ),
.I2(CLBLL_L_X42Y96_SLICE_X69Y96_B5Q),
.I3(CLBLL_L_X42Y118_SLICE_X69Y118_C5Q),
.I4(CLBLL_L_X42Y118_SLICE_X69Y118_BQ),
.I5(CLBLL_L_X42Y118_SLICE_X69Y118_AQ),
.O5(CLBLL_L_X42Y96_SLICE_X69Y96_DO5),
.O6(CLBLL_L_X42Y96_SLICE_X69Y96_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccf0f0ff00aaaa)
  ) CLBLL_L_X42Y96_SLICE_X69Y96_CLUT (
.I0(CLBLL_L_X42Y118_SLICE_X69Y118_B5Q),
.I1(CLBLL_L_X42Y118_SLICE_X69Y118_A5Q),
.I2(CLBLL_L_X42Y118_SLICE_X69Y118_CQ),
.I3(CLBLL_L_X42Y118_SLICE_X69Y118_D5Q),
.I4(CLBLL_L_X42Y96_SLICE_X69Y96_BQ),
.I5(CLBLL_L_X42Y96_SLICE_X69Y96_B5Q),
.O5(CLBLL_L_X42Y96_SLICE_X69Y96_CO5),
.O6(CLBLL_L_X42Y96_SLICE_X69Y96_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0fcccccccc)
  ) CLBLL_L_X42Y96_SLICE_X69Y96_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y96_SLICE_X69Y96_AO6),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y96_SLICE_X69Y96_BO5),
.O6(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcaaaeaaa0aaa2aaa)
  ) CLBLL_L_X42Y96_SLICE_X69Y96_ALUT (
.I0(CLBLL_L_X42Y96_SLICE_X69Y96_BQ),
.I1(CLBLL_L_X42Y112_SLICE_X69Y112_C5Q),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(CLBLL_L_X42Y71_SLICE_X68Y71_BQ),
.I4(CLBLL_L_X42Y112_SLICE_X69Y112_DQ),
.I5(CLBLL_L_X42Y43_SLICE_X68Y43_C_XOR),
.O5(CLBLL_L_X42Y96_SLICE_X69Y96_AO5),
.O6(CLBLL_L_X42Y96_SLICE_X69Y96_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y97_SLICE_X68Y97_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y97_SLICE_X68Y97_AO6),
.Q(CLBLL_L_X42Y97_SLICE_X68Y97_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y97_SLICE_X68Y97_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(1'b1),
.D(CLBLL_L_X42Y97_SLICE_X68Y97_AO5),
.Q(CLBLL_L_X42Y97_SLICE_X68Y97_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000002)
  ) CLBLL_L_X42Y97_SLICE_X68Y97_DLUT (
.I0(CLBLL_L_X42Y97_SLICE_X68Y97_BO5),
.I1(CLBLL_L_X42Y93_SLICE_X68Y93_BQ),
.I2(CLBLL_L_X42Y93_SLICE_X68Y93_DQ),
.I3(CLBLL_L_X42Y104_SLICE_X69Y104_CQ),
.I4(CLBLL_L_X42Y93_SLICE_X68Y93_CQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y97_SLICE_X68Y97_DO5),
.O6(CLBLL_L_X42Y97_SLICE_X68Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h1000a0a00010a0a0)
  ) CLBLL_L_X42Y97_SLICE_X68Y97_CLUT (
.I0(CLBLL_L_X42Y113_SLICE_X68Y113_D5Q),
.I1(CLBLL_L_X42Y92_SLICE_X69Y92_B5Q),
.I2(CLBLL_L_X42Y97_SLICE_X68Y97_DO5),
.I3(CLBLL_L_X42Y95_SLICE_X68Y95_D5Q),
.I4(CLBLL_L_X42Y93_SLICE_X68Y93_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X42Y97_SLICE_X68Y97_CO5),
.O6(CLBLL_L_X42Y97_SLICE_X68Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'ha0a0a0a000330033)
  ) CLBLL_L_X42Y97_SLICE_X68Y97_BLUT (
.I0(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I1(CLBLL_L_X42Y104_SLICE_X69Y104_BQ),
.I2(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I3(CLBLL_L_X42Y104_SLICE_X69Y104_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y97_SLICE_X68Y97_BO5),
.O6(CLBLL_L_X42Y97_SLICE_X68Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000bf3f8000)
  ) CLBLL_L_X42Y97_SLICE_X68Y97_ALUT (
.I0(CLBLL_L_X42Y93_SLICE_X68Y93_B_XOR),
.I1(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(CLBLL_L_X42Y96_SLICE_X68Y96_AO5),
.I4(CLBLL_L_X42Y97_SLICE_X68Y97_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y97_SLICE_X68Y97_AO5),
.O6(CLBLL_L_X42Y97_SLICE_X68Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y97_SLICE_X69Y97_C5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X68Y97_CO5),
.D(CLBLL_L_X42Y97_SLICE_X69Y97_CO5),
.Q(CLBLL_L_X42Y97_SLICE_X69Y97_C5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hd00d000000000000)
  ) CLBLL_L_X42Y97_SLICE_X69Y97_DLUT (
.I0(BRAM_L_X44Y95_RAMB18_X2Y38_DO7),
.I1(CLBLL_L_X42Y95_SLICE_X69Y95_D5Q),
.I2(BRAM_L_X44Y95_RAMB18_X2Y38_DO2),
.I3(CLBLL_L_X42Y95_SLICE_X69Y95_AQ),
.I4(CLBLL_L_X42Y97_SLICE_X69Y97_AO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y97_SLICE_X69Y97_DO5),
.O6(CLBLL_L_X42Y97_SLICE_X69Y97_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100010055550000)
  ) CLBLL_L_X42Y97_SLICE_X69Y97_CLUT (
.I0(CLBLL_L_X42Y97_SLICE_X69Y97_BO5),
.I1(CLBLL_L_X42Y92_SLICE_X69Y92_B5Q),
.I2(CLBLL_L_X42Y95_SLICE_X68Y95_D5Q),
.I3(CLBLL_L_X42Y97_SLICE_X68Y97_BO6),
.I4(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y97_SLICE_X69Y97_CO5),
.O6(CLBLL_L_X42Y97_SLICE_X69Y97_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000088002200)
  ) CLBLL_L_X42Y97_SLICE_X69Y97_BLUT (
.I0(CLBLL_L_X42Y97_SLICE_X69Y97_DO6),
.I1(BRAM_L_X44Y95_RAMB18_X2Y38_DO5),
.I2(1'b1),
.I3(CLBLL_L_X42Y93_SLICE_X69Y93_CO5),
.I4(CLBLL_L_X42Y91_SLICE_X69Y91_D5Q),
.I5(1'b1),
.O5(CLBLL_L_X42Y97_SLICE_X69Y97_BO5),
.O6(CLBLL_L_X42Y97_SLICE_X69Y97_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0300000301000001)
  ) CLBLL_L_X42Y97_SLICE_X69Y97_ALUT (
.I0(BRAM_L_X44Y95_RAMB18_X2Y38_DO4),
.I1(BRAM_L_X44Y95_RAMB18_X2Y38_DO10),
.I2(BRAM_L_X44Y95_RAMB18_X2Y38_DO9),
.I3(BRAM_L_X44Y95_RAMB18_X2Y38_DOP0),
.I4(CLBLL_L_X42Y95_SLICE_X69Y95_CQ),
.I5(CLBLL_L_X42Y92_SLICE_X69Y92_AQ),
.O5(CLBLL_L_X42Y97_SLICE_X69Y97_AO5),
.O6(CLBLL_L_X42Y97_SLICE_X69Y97_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y98_SLICE_X68Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y98_SLICE_X68Y98_DO5),
.O6(CLBLL_L_X42Y98_SLICE_X68Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y98_SLICE_X68Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y98_SLICE_X68Y98_CO5),
.O6(CLBLL_L_X42Y98_SLICE_X68Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y98_SLICE_X68Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y98_SLICE_X68Y98_BO5),
.O6(CLBLL_L_X42Y98_SLICE_X68Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y98_SLICE_X68Y98_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y98_SLICE_X68Y98_AO5),
.O6(CLBLL_L_X42Y98_SLICE_X68Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y98_SLICE_X69Y98_D5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(BRAM_L_X44Y95_RAMB18_X2Y38_DO6),
.Q(CLBLL_L_X42Y98_SLICE_X69Y98_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y98_SLICE_X69Y98_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(BRAM_L_X44Y95_RAMB18_X2Y38_DO8),
.Q(CLBLL_L_X42Y98_SLICE_X69Y98_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y98_SLICE_X69Y98_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y98_SLICE_X69Y98_DO5),
.O6(CLBLL_L_X42Y98_SLICE_X69Y98_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y98_SLICE_X69Y98_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y98_SLICE_X69Y98_CO5),
.O6(CLBLL_L_X42Y98_SLICE_X69Y98_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y98_SLICE_X69Y98_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y98_SLICE_X69Y98_BO5),
.O6(CLBLL_L_X42Y98_SLICE_X69Y98_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y98_SLICE_X69Y98_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y98_SLICE_X69Y98_AO5),
.O6(CLBLL_L_X42Y98_SLICE_X69Y98_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y101_SLICE_X68Y101_A5_FDSE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y71_SLICE_X68Y71_BQ),
.D(CLBLL_L_X42Y101_SLICE_X68Y101_AO5),
.Q(CLBLL_L_X42Y101_SLICE_X68Y101_A5Q),
.S(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y101_SLICE_X68Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y101_SLICE_X68Y101_DO5),
.O6(CLBLL_L_X42Y101_SLICE_X68Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y101_SLICE_X68Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y101_SLICE_X68Y101_CO5),
.O6(CLBLL_L_X42Y101_SLICE_X68Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y101_SLICE_X68Y101_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y101_SLICE_X68Y101_BO5),
.O6(CLBLL_L_X42Y101_SLICE_X68Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000e020ef2f)
  ) CLBLL_L_X42Y101_SLICE_X68Y101_ALUT (
.I0(CLBLL_L_X42Y96_SLICE_X69Y96_DO6),
.I1(CLBLL_L_X42Y110_SLICE_X69Y110_C5Q),
.I2(CLBLL_L_X42Y112_SLICE_X69Y112_C5Q),
.I3(CLBLL_L_X42Y96_SLICE_X69Y96_CO6),
.I4(CLBLL_L_X42Y112_SLICE_X69Y112_DQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y101_SLICE_X68Y101_AO5),
.O6(CLBLL_L_X42Y101_SLICE_X68Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y101_SLICE_X69Y101_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y101_SLICE_X69Y101_AO5),
.Q(CLBLL_L_X42Y101_SLICE_X69Y101_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y101_SLICE_X69Y101_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y101_SLICE_X69Y101_CO5),
.Q(CLBLL_L_X42Y101_SLICE_X69Y101_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y101_SLICE_X69Y101_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y95_SLICE_X69Y95_AQ),
.Q(CLBLL_L_X42Y101_SLICE_X69Y101_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y101_SLICE_X69Y101_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y95_SLICE_X69Y95_D5Q),
.Q(CLBLL_L_X42Y101_SLICE_X69Y101_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y101_SLICE_X69Y101_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y95_SLICE_X69Y95_CQ),
.Q(CLBLL_L_X42Y101_SLICE_X69Y101_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y101_SLICE_X69Y101_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y91_SLICE_X69Y91_D5Q),
.Q(CLBLL_L_X42Y101_SLICE_X69Y101_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h15153f3f00000000)
  ) CLBLL_L_X42Y101_SLICE_X69Y101_DLUT (
.I0(CLBLL_L_X42Y107_SLICE_X68Y107_BO5),
.I1(CLBLL_L_X42Y106_SLICE_X69Y106_CO5),
.I2(CLBLL_L_X42Y68_SLICE_X68Y68_A5Q),
.I3(1'b1),
.I4(CLBLM_R_X41Y95_SLICE_X67Y95_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y101_SLICE_X69Y101_DO5),
.O6(CLBLL_L_X42Y101_SLICE_X69Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLL_L_X42Y101_SLICE_X69Y101_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X42Y91_SLICE_X69Y91_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y101_SLICE_X69Y101_CO5),
.O6(CLBLL_L_X42Y101_SLICE_X69Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000033ff33)
  ) CLBLL_L_X42Y101_SLICE_X69Y101_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X41Y111_SLICE_X66Y111_BQ),
.I2(1'b1),
.I3(CLBLL_L_X42Y106_SLICE_X69Y106_CO5),
.I4(CLBLL_L_X42Y68_SLICE_X68Y68_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X42Y101_SLICE_X69Y101_BO5),
.O6(CLBLL_L_X42Y101_SLICE_X69Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaaaaaa)
  ) CLBLL_L_X42Y101_SLICE_X69Y101_ALUT (
.I0(BRAM_L_X44Y95_RAMB18_X2Y38_DO11),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y101_SLICE_X69Y101_AO5),
.O6(CLBLL_L_X42Y101_SLICE_X69Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y102_SLICE_X68Y102_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y102_SLICE_X68Y102_DO5),
.D(CLBLL_L_X42Y102_SLICE_X68Y102_BO6),
.Q(CLBLL_L_X42Y102_SLICE_X68Y102_BQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000333300a200a2)
  ) CLBLL_L_X42Y102_SLICE_X68Y102_DLUT (
.I0(CLBLL_L_X42Y102_SLICE_X68Y102_CO5),
.I1(CLBLL_L_X42Y109_SLICE_X69Y109_CO6),
.I2(CLBLL_L_X42Y103_SLICE_X68Y103_CO6),
.I3(CLBLM_R_X41Y115_SLICE_X66Y115_DO6),
.I4(CLBLM_R_X41Y107_SLICE_X66Y107_AO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y102_SLICE_X68Y102_DO5),
.O6(CLBLL_L_X42Y102_SLICE_X68Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc0000f055ff)
  ) CLBLL_L_X42Y102_SLICE_X68Y102_CLUT (
.I0(CLBLM_R_X41Y102_SLICE_X66Y102_BO5),
.I1(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I2(CLBLM_R_X41Y102_SLICE_X66Y102_CO6),
.I3(CLBLM_R_X41Y109_SLICE_X67Y109_CO6),
.I4(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y102_SLICE_X68Y102_CO5),
.O6(CLBLL_L_X42Y102_SLICE_X68Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcf05cf050000cccc)
  ) CLBLL_L_X42Y102_SLICE_X68Y102_BLUT (
.I0(CLBLL_L_X42Y102_SLICE_X68Y102_AO6),
.I1(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I2(CLBLM_R_X41Y102_SLICE_X66Y102_CO6),
.I3(CLBLL_L_X42Y110_SLICE_X69Y110_BO6),
.I4(CLBLM_R_X41Y107_SLICE_X67Y107_D5Q),
.I5(1'b1),
.O5(CLBLL_L_X42Y102_SLICE_X68Y102_BO5),
.O6(CLBLL_L_X42Y102_SLICE_X68Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ff000000550000)
  ) CLBLL_L_X42Y102_SLICE_X68Y102_ALUT (
.I0(CLBLL_L_X42Y102_SLICE_X68Y102_DO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X42Y103_SLICE_X69Y103_B_XOR),
.I4(CLBLL_L_X42Y103_SLICE_X69Y103_AO5),
.I5(1'b1),
.O5(CLBLL_L_X42Y102_SLICE_X68Y102_AO5),
.O6(CLBLL_L_X42Y102_SLICE_X68Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y102_SLICE_X69Y102_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y102_SLICE_X69Y102_AO5),
.Q(CLBLL_L_X42Y102_SLICE_X69Y102_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y102_SLICE_X69Y102_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y102_SLICE_X69Y102_CO5),
.Q(CLBLL_L_X42Y102_SLICE_X69Y102_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y102_SLICE_X69Y102_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y102_SLICE_X69Y102_DO5),
.Q(CLBLL_L_X42Y102_SLICE_X69Y102_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y102_SLICE_X69Y102_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y112_SLICE_X68Y112_D5Q),
.Q(CLBLL_L_X42Y102_SLICE_X69Y102_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y102_SLICE_X69Y102_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y113_SLICE_X69Y113_A5Q),
.Q(CLBLL_L_X42Y102_SLICE_X69Y102_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y102_SLICE_X69Y102_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y101_SLICE_X69Y101_D5Q),
.Q(CLBLL_L_X42Y102_SLICE_X69Y102_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaaaaaa)
  ) CLBLL_L_X42Y102_SLICE_X69Y102_DLUT (
.I0(CLBLL_L_X42Y111_SLICE_X68Y111_B5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y102_SLICE_X69Y102_DO5),
.O6(CLBLL_L_X42Y102_SLICE_X69Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLL_L_X42Y102_SLICE_X69Y102_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X42Y112_SLICE_X68Y112_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y102_SLICE_X69Y102_CO5),
.O6(CLBLL_L_X42Y102_SLICE_X69Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000ff2727)
  ) CLBLL_L_X42Y102_SLICE_X69Y102_BLUT (
.I0(CLBLL_L_X42Y106_SLICE_X69Y106_CO5),
.I1(CLBLL_L_X42Y102_SLICE_X69Y102_D5Q),
.I2(CLBLL_L_X42Y102_SLICE_X69Y102_DQ),
.I3(CLBLL_L_X42Y102_SLICE_X69Y102_A5Q),
.I4(CLBLL_L_X42Y102_SLICE_X68Y102_CO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y102_SLICE_X69Y102_BO5),
.O6(CLBLL_L_X42Y102_SLICE_X69Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff0000)
  ) CLBLL_L_X42Y102_SLICE_X69Y102_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X42Y112_SLICE_X68Y112_DQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y102_SLICE_X69Y102_AO5),
.O6(CLBLL_L_X42Y102_SLICE_X69Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y103_SLICE_X68Y103_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y103_SLICE_X68Y103_DO5),
.D(CLBLL_L_X42Y104_SLICE_X69Y104_BO5),
.Q(CLBLL_L_X42Y103_SLICE_X68Y103_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y103_SLICE_X68Y103_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y103_SLICE_X68Y103_DO5),
.D(CLBLL_L_X42Y104_SLICE_X69Y104_CO5),
.Q(CLBLL_L_X42Y103_SLICE_X68Y103_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y103_SLICE_X68Y103_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y103_SLICE_X68Y103_DO5),
.D(CLBLL_L_X42Y104_SLICE_X69Y104_DO5),
.Q(CLBLL_L_X42Y103_SLICE_X68Y103_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000005000)
  ) CLBLL_L_X42Y103_SLICE_X68Y103_DLUT (
.I0(CLBLL_L_X42Y109_SLICE_X69Y109_BO5),
.I1(1'b1),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(CLBLL_L_X42Y103_SLICE_X68Y103_CO5),
.I4(CLBLM_R_X41Y109_SLICE_X66Y109_BO5),
.I5(1'b1),
.O5(CLBLL_L_X42Y103_SLICE_X68Y103_DO5),
.O6(CLBLL_L_X42Y103_SLICE_X68Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000333300aaccff)
  ) CLBLL_L_X42Y103_SLICE_X68Y103_CLUT (
.I0(CLBLL_L_X42Y102_SLICE_X68Y102_DO6),
.I1(CLBLL_L_X42Y102_SLICE_X68Y102_AO6),
.I2(1'b1),
.I3(CLBLM_R_X41Y108_SLICE_X67Y108_BO6),
.I4(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y103_SLICE_X68Y103_CO5),
.O6(CLBLL_L_X42Y103_SLICE_X68Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000050005)
  ) CLBLL_L_X42Y103_SLICE_X68Y103_BLUT (
.I0(CLBLL_L_X42Y103_SLICE_X68Y103_CQ),
.I1(1'b1),
.I2(CLBLL_L_X42Y103_SLICE_X68Y103_DQ),
.I3(CLBLL_L_X42Y103_SLICE_X68Y103_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.O6(CLBLL_L_X42Y103_SLICE_X68Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h05000d0000000800)
  ) CLBLL_L_X42Y103_SLICE_X68Y103_ALUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I1(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I2(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I3(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I4(CLBLM_R_X41Y106_SLICE_X66Y106_CO6),
.I5(CLBLM_R_X41Y105_SLICE_X66Y105_CO6),
.O5(CLBLL_L_X42Y103_SLICE_X68Y103_AO5),
.O6(CLBLL_L_X42Y103_SLICE_X68Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y103_SLICE_X69Y103_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y103_SLICE_X68Y103_DO5),
.D(CLBLL_L_X42Y103_SLICE_X69Y103_BO5),
.Q(CLBLL_L_X42Y103_SLICE_X69Y103_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X42Y103_SLICE_X69Y103_CARRY4 (
.CI(1'b0),
.CO({CLBLL_L_X42Y103_SLICE_X69Y103_D_CY, CLBLL_L_X42Y103_SLICE_X69Y103_C_CY, CLBLL_L_X42Y103_SLICE_X69Y103_B_CY, CLBLL_L_X42Y103_SLICE_X69Y103_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({CLBLL_L_X42Y103_SLICE_X69Y103_D_XOR, CLBLL_L_X42Y103_SLICE_X69Y103_C_XOR, CLBLL_L_X42Y103_SLICE_X69Y103_B_XOR, CLBLL_L_X42Y103_SLICE_X69Y103_A_XOR}),
.S({CLBLL_L_X42Y103_SLICE_X69Y103_DO6, CLBLL_L_X42Y103_SLICE_X69Y103_CO6, CLBLL_L_X42Y103_SLICE_X69Y103_BO6, CLBLL_L_X42Y103_SLICE_X69Y103_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000000000)
  ) CLBLL_L_X42Y103_SLICE_X69Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X42Y103_SLICE_X68Y103_CQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y103_SLICE_X69Y103_DO5),
.O6(CLBLL_L_X42Y103_SLICE_X69Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLL_L_X42Y103_SLICE_X69Y103_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X42Y103_SLICE_X68Y103_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y103_SLICE_X69Y103_CO5),
.O6(CLBLL_L_X42Y103_SLICE_X69Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0fcccf000)
  ) CLBLL_L_X42Y103_SLICE_X69Y103_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y103_SLICE_X69Y103_B_XOR),
.I2(CLBLL_L_X42Y103_SLICE_X69Y103_BQ),
.I3(CLBLL_L_X42Y110_SLICE_X68Y110_BO5),
.I4(CLBLM_R_X41Y108_SLICE_X67Y108_BO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y103_SLICE_X69Y103_BO5),
.O6(CLBLL_L_X42Y103_SLICE_X69Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000110011)
  ) CLBLL_L_X42Y103_SLICE_X69Y103_ALUT (
.I0(CLBLL_L_X42Y103_SLICE_X69Y103_C_XOR),
.I1(CLBLL_L_X42Y104_SLICE_X69Y104_A_XOR),
.I2(CLBLL_L_X42Y104_SLICE_X68Y104_DO5),
.I3(CLBLL_L_X42Y103_SLICE_X69Y103_D_XOR),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y103_SLICE_X69Y103_AO5),
.O6(CLBLL_L_X42Y103_SLICE_X69Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y104_SLICE_X68Y104_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y103_SLICE_X68Y103_DO5),
.D(CLBLL_L_X42Y108_SLICE_X69Y108_CO5),
.Q(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccffcc000f0f0f0f)
  ) CLBLL_L_X42Y104_SLICE_X68Y104_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y105_SLICE_X69Y105_BO6),
.I2(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.I3(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I4(CLBLM_R_X41Y106_SLICE_X67Y106_BO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y104_SLICE_X68Y104_DO5),
.O6(CLBLL_L_X42Y104_SLICE_X68Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h54040000feae0000)
  ) CLBLL_L_X42Y104_SLICE_X68Y104_CLUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I1(CLBLM_R_X41Y106_SLICE_X67Y106_BO6),
.I2(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I3(CLBLL_L_X42Y105_SLICE_X69Y105_BO6),
.I4(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.I5(CLBLL_L_X42Y104_SLICE_X68Y104_AO6),
.O5(CLBLL_L_X42Y104_SLICE_X68Y104_CO5),
.O6(CLBLL_L_X42Y104_SLICE_X68Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5000202050007070)
  ) CLBLL_L_X42Y104_SLICE_X68Y104_BLUT (
.I0(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.I1(CLBLL_L_X42Y104_SLICE_X68Y104_AO6),
.I2(CLBLM_R_X41Y107_SLICE_X67Y107_BO6),
.I3(CLBLL_L_X42Y104_SLICE_X68Y104_DO6),
.I4(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I5(CLBLM_R_X41Y105_SLICE_X66Y105_AO6),
.O5(CLBLL_L_X42Y104_SLICE_X68Y104_BO5),
.O6(CLBLL_L_X42Y104_SLICE_X68Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5515ffbf1115bbbf)
  ) CLBLL_L_X42Y104_SLICE_X68Y104_ALUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I1(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I2(CLBLL_L_X42Y106_SLICE_X68Y106_DO5),
.I3(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I4(CLBLL_L_X42Y105_SLICE_X68Y105_BO5),
.I5(CLBLL_L_X42Y101_SLICE_X69Y101_DO6),
.O5(CLBLL_L_X42Y104_SLICE_X68Y104_AO5),
.O6(CLBLL_L_X42Y104_SLICE_X68Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y104_SLICE_X69Y104_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.D(1'b0),
.Q(CLBLL_L_X42Y104_SLICE_X69Y104_AQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y104_SLICE_X69Y104_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.D(1'b0),
.Q(CLBLL_L_X42Y104_SLICE_X69Y104_BQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y104_SLICE_X69Y104_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X68Y97_CO6),
.D(1'b0),
.Q(CLBLL_L_X42Y104_SLICE_X69Y104_CQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X42Y104_SLICE_X69Y104_CARRY4 (
.CI(CLBLL_L_X42Y103_SLICE_X69Y103_COUT),
.CO({CLBLL_L_X42Y104_SLICE_X69Y104_COUT, CLBLL_L_X42Y104_SLICE_X69Y104_C_CY, CLBLL_L_X42Y104_SLICE_X69Y104_B_CY, CLBLL_L_X42Y104_SLICE_X69Y104_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLL_L_X42Y104_SLICE_X69Y104_D_XOR, CLBLL_L_X42Y104_SLICE_X69Y104_C_XOR, CLBLL_L_X42Y104_SLICE_X69Y104_B_XOR, CLBLL_L_X42Y104_SLICE_X69Y104_A_XOR}),
.S({CLBLL_L_X42Y104_SLICE_X69Y104_DO6, CLBLL_L_X42Y104_SLICE_X69Y104_CO6, CLBLL_L_X42Y104_SLICE_X69Y104_BO6, CLBLL_L_X42Y104_SLICE_X69Y104_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00f8f88888)
  ) CLBLL_L_X42Y104_SLICE_X69Y104_DLUT (
.I0(CLBLL_L_X42Y103_SLICE_X68Y103_DQ),
.I1(CLBLL_L_X42Y110_SLICE_X68Y110_BO5),
.I2(CLBLM_R_X41Y108_SLICE_X67Y108_BO6),
.I3(1'b0),
.I4(CLBLL_L_X42Y103_SLICE_X69Y103_C_XOR),
.I5(1'b1),
.O5(CLBLL_L_X42Y104_SLICE_X69Y104_DO5),
.O6(CLBLL_L_X42Y104_SLICE_X69Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff888888)
  ) CLBLL_L_X42Y104_SLICE_X69Y104_CLUT (
.I0(CLBLL_L_X42Y103_SLICE_X69Y103_D_XOR),
.I1(CLBLM_R_X41Y108_SLICE_X67Y108_BO6),
.I2(1'b0),
.I3(CLBLL_L_X42Y110_SLICE_X68Y110_BO5),
.I4(CLBLL_L_X42Y103_SLICE_X68Y103_CQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y104_SLICE_X69Y104_CO5),
.O6(CLBLL_L_X42Y104_SLICE_X69Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f888f888)
  ) CLBLL_L_X42Y104_SLICE_X69Y104_BLUT (
.I0(CLBLM_R_X41Y108_SLICE_X67Y108_BO6),
.I1(CLBLL_L_X42Y104_SLICE_X69Y104_A_XOR),
.I2(CLBLL_L_X42Y103_SLICE_X68Y103_BQ),
.I3(CLBLL_L_X42Y110_SLICE_X68Y110_BO5),
.I4(1'b0),
.I5(1'b1),
.O5(CLBLL_L_X42Y104_SLICE_X69Y104_BO5),
.O6(CLBLL_L_X42Y104_SLICE_X69Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLL_L_X42Y104_SLICE_X69Y104_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y103_SLICE_X68Y103_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y104_SLICE_X69Y104_AO5),
.O6(CLBLL_L_X42Y104_SLICE_X69Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y105_SLICE_X68Y105_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y92_SLICE_X68Y92_CQ),
.Q(CLBLL_L_X42Y105_SLICE_X68Y105_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'ha2aaf7ff02aa57ff)
  ) CLBLL_L_X42Y105_SLICE_X68Y105_DLUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I1(CLBLL_L_X42Y106_SLICE_X68Y106_DO5),
.I2(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I3(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I4(CLBLL_L_X42Y105_SLICE_X69Y105_BO6),
.I5(CLBLL_L_X42Y101_SLICE_X69Y101_DO6),
.O5(CLBLL_L_X42Y105_SLICE_X68Y105_DO5),
.O6(CLBLL_L_X42Y105_SLICE_X68Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf3f3c0c022222222)
  ) CLBLL_L_X42Y105_SLICE_X68Y105_CLUT (
.I0(CLBLL_L_X42Y105_SLICE_X68Y105_BO5),
.I1(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I2(CLBLM_R_X41Y106_SLICE_X67Y106_BO6),
.I3(1'b1),
.I4(CLBLM_R_X41Y106_SLICE_X66Y106_AO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y105_SLICE_X68Y105_CO5),
.O6(CLBLL_L_X42Y105_SLICE_X68Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000e0a0c000)
  ) CLBLL_L_X42Y105_SLICE_X68Y105_BLUT (
.I0(CLBLL_L_X42Y105_SLICE_X68Y105_CQ),
.I1(CLBLM_R_X41Y114_SLICE_X67Y114_DQ),
.I2(CLBLL_L_X42Y106_SLICE_X69Y106_DO5),
.I3(CLBLL_L_X42Y107_SLICE_X68Y107_BO5),
.I4(CLBLL_L_X42Y106_SLICE_X69Y106_CO5),
.I5(1'b1),
.O5(CLBLL_L_X42Y105_SLICE_X68Y105_BO5),
.O6(CLBLL_L_X42Y105_SLICE_X68Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h45004f0040004a00)
  ) CLBLL_L_X42Y105_SLICE_X68Y105_ALUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I1(CLBLL_L_X42Y105_SLICE_X68Y105_CO5),
.I2(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.I3(CLBLM_R_X41Y107_SLICE_X67Y107_BO6),
.I4(CLBLL_L_X42Y105_SLICE_X68Y105_DO6),
.I5(CLBLL_L_X42Y105_SLICE_X68Y105_CO6),
.O5(CLBLL_L_X42Y105_SLICE_X68Y105_AO5),
.O6(CLBLL_L_X42Y105_SLICE_X68Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y105_SLICE_X69Y105_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y105_SLICE_X69Y105_AO5),
.Q(CLBLL_L_X42Y105_SLICE_X69Y105_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y105_SLICE_X69Y105_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y101_SLICE_X69Y101_AQ),
.Q(CLBLL_L_X42Y105_SLICE_X69Y105_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000c0a0c000)
  ) CLBLL_L_X42Y105_SLICE_X69Y105_DLUT (
.I0(CLBLM_R_X41Y108_SLICE_X67Y108_CO6),
.I1(CLBLM_R_X41Y95_SLICE_X67Y95_DQ),
.I2(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I3(CLBLL_L_X42Y106_SLICE_X69Y106_CO6),
.I4(CLBLL_L_X42Y111_SLICE_X69Y111_D5Q),
.I5(1'b1),
.O5(CLBLL_L_X42Y105_SLICE_X69Y105_DO5),
.O6(CLBLL_L_X42Y105_SLICE_X69Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cac00000)
  ) CLBLL_L_X42Y105_SLICE_X69Y105_CLUT (
.I0(CLBLL_L_X42Y105_SLICE_X69Y105_A5Q),
.I1(CLBLM_R_X41Y95_SLICE_X67Y95_CQ),
.I2(CLBLL_L_X42Y106_SLICE_X69Y106_CO6),
.I3(CLBLM_R_X41Y108_SLICE_X67Y108_CO6),
.I4(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y105_SLICE_X69Y105_CO5),
.O6(CLBLL_L_X42Y105_SLICE_X69Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf5a00000d8d80000)
  ) CLBLL_L_X42Y105_SLICE_X69Y105_BLUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I1(CLBLL_L_X42Y106_SLICE_X68Y106_DO5),
.I2(CLBLL_L_X42Y105_SLICE_X69Y105_CO5),
.I3(CLBLL_L_X42Y105_SLICE_X69Y105_DO5),
.I4(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I5(1'b1),
.O5(CLBLL_L_X42Y105_SLICE_X69Y105_BO5),
.O6(CLBLL_L_X42Y105_SLICE_X69Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f0f0f0f0)
  ) CLBLL_L_X42Y105_SLICE_X69Y105_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y101_SLICE_X69Y101_A5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y105_SLICE_X69Y105_AO5),
.O6(CLBLL_L_X42Y105_SLICE_X69Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y106_SLICE_X68Y106_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y106_SLICE_X68Y106_AO5),
.Q(CLBLL_L_X42Y106_SLICE_X68Y106_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y106_SLICE_X68Y106_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y113_SLICE_X69Y113_CQ),
.Q(CLBLL_L_X42Y106_SLICE_X68Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000e4a00000)
  ) CLBLL_L_X42Y106_SLICE_X68Y106_DLUT (
.I0(CLBLL_L_X42Y106_SLICE_X69Y106_CO6),
.I1(CLBLL_L_X42Y107_SLICE_X69Y107_C5Q),
.I2(CLBLM_R_X41Y95_SLICE_X67Y95_AQ),
.I3(CLBLM_R_X41Y108_SLICE_X67Y108_CO6),
.I4(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y106_SLICE_X68Y106_DO5),
.O6(CLBLL_L_X42Y106_SLICE_X68Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000135f5f5f)
  ) CLBLL_L_X42Y106_SLICE_X68Y106_CLUT (
.I0(CLBLL_L_X42Y106_SLICE_X69Y106_CO5),
.I1(CLBLM_R_X41Y114_SLICE_X67Y114_DQ),
.I2(CLBLL_L_X42Y105_SLICE_X68Y105_CQ),
.I3(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I4(CLBLM_R_X41Y107_SLICE_X66Y107_AO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y106_SLICE_X68Y106_CO5),
.O6(CLBLL_L_X42Y106_SLICE_X68Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000078f070f)
  ) CLBLL_L_X42Y106_SLICE_X68Y106_BLUT (
.I0(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I1(CLBLL_L_X42Y109_SLICE_X69Y109_BO6),
.I2(CLBLL_L_X42Y106_SLICE_X68Y106_AQ),
.I3(CLBLL_L_X42Y106_SLICE_X68Y106_A5Q),
.I4(CLBLL_L_X42Y108_SLICE_X68Y108_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X42Y106_SLICE_X68Y106_BO5),
.O6(CLBLL_L_X42Y106_SLICE_X68Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff0000)
  ) CLBLL_L_X42Y106_SLICE_X68Y106_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X42Y98_SLICE_X69Y98_D5Q),
.I5(1'b1),
.O5(CLBLL_L_X42Y106_SLICE_X68Y106_AO5),
.O6(CLBLL_L_X42Y106_SLICE_X68Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y106_SLICE_X69Y106_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y80_SLICE_X69Y80_B5Q),
.Q(CLBLL_L_X42Y106_SLICE_X69Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaccaacc0f0f0000)
  ) CLBLL_L_X42Y106_SLICE_X69Y106_DLUT (
.I0(CLBLL_L_X42Y106_SLICE_X69Y106_CQ),
.I1(CLBLL_L_X42Y68_SLICE_X68Y68_CQ),
.I2(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I3(CLBLL_L_X42Y106_SLICE_X69Y106_CO5),
.I4(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I5(1'b1),
.O5(CLBLL_L_X42Y106_SLICE_X69Y106_DO5),
.O6(CLBLL_L_X42Y106_SLICE_X69Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000330000220000)
  ) CLBLL_L_X42Y106_SLICE_X69Y106_CLUT (
.I0(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I1(CLBLM_R_X41Y102_SLICE_X67Y102_C5Q),
.I2(1'b1),
.I3(CLBLL_L_X42Y109_SLICE_X69Y109_DQ),
.I4(CLBLL_L_X42Y108_SLICE_X68Y108_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X42Y106_SLICE_X69Y106_CO5),
.O6(CLBLL_L_X42Y106_SLICE_X69Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000011151515)
  ) CLBLL_L_X42Y106_SLICE_X69Y106_BLUT (
.I0(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.I1(CLBLM_R_X41Y105_SLICE_X67Y105_CO6),
.I2(CLBLL_L_X42Y106_SLICE_X69Y106_AO6),
.I3(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I4(CLBLL_L_X42Y107_SLICE_X68Y107_CO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y106_SLICE_X69Y106_BO5),
.O6(CLBLL_L_X42Y106_SLICE_X69Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa008a8aaa008080)
  ) CLBLL_L_X42Y106_SLICE_X69Y106_ALUT (
.I0(CLBLL_L_X42Y106_SLICE_X69Y106_DO5),
.I1(CLBLL_L_X42Y108_SLICE_X69Y108_AQ),
.I2(CLBLM_R_X41Y108_SLICE_X66Y108_CO6),
.I3(CLBLM_R_X41Y100_SLICE_X67Y100_AQ),
.I4(CLBLL_L_X42Y107_SLICE_X68Y107_BO5),
.I5(CLBLL_L_X42Y106_SLICE_X69Y106_DO6),
.O5(CLBLL_L_X42Y106_SLICE_X69Y106_AO5),
.O6(CLBLL_L_X42Y106_SLICE_X69Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y107_SLICE_X68Y107_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y101_SLICE_X69Y101_C5Q),
.Q(CLBLL_L_X42Y107_SLICE_X68Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000f0f000ff407f)
  ) CLBLL_L_X42Y107_SLICE_X68Y107_DLUT (
.I0(CLBLL_L_X42Y68_SLICE_X68Y68_DQ),
.I1(CLBLM_R_X41Y108_SLICE_X67Y108_BO6),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(CLBLL_L_X42Y107_SLICE_X68Y107_BQ),
.I4(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y107_SLICE_X68Y107_DO5),
.O6(CLBLL_L_X42Y107_SLICE_X68Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hb0808080b0b080b0)
  ) CLBLL_L_X42Y107_SLICE_X68Y107_CLUT (
.I0(CLBLM_R_X41Y100_SLICE_X67Y100_D5Q),
.I1(CLBLL_L_X42Y107_SLICE_X68Y107_BO5),
.I2(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I3(CLBLM_R_X41Y108_SLICE_X66Y108_CO6),
.I4(CLBLL_L_X42Y107_SLICE_X69Y107_AQ),
.I5(CLBLL_L_X42Y101_SLICE_X69Y101_BO5),
.O5(CLBLL_L_X42Y107_SLICE_X68Y107_CO5),
.O6(CLBLL_L_X42Y107_SLICE_X68Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf7f7000088888888)
  ) CLBLL_L_X42Y107_SLICE_X68Y107_BLUT (
.I0(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I1(CLBLM_R_X41Y107_SLICE_X66Y107_AO6),
.I2(CLBLM_R_X41Y106_SLICE_X67Y106_C5Q),
.I3(1'b1),
.I4(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I5(1'b1),
.O5(CLBLL_L_X42Y107_SLICE_X68Y107_BO5),
.O6(CLBLL_L_X42Y107_SLICE_X68Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcc00cc008c8c0404)
  ) CLBLL_L_X42Y107_SLICE_X68Y107_ALUT (
.I0(CLBLM_R_X41Y108_SLICE_X66Y108_CO6),
.I1(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I2(CLBLL_L_X42Y107_SLICE_X68Y107_DO5),
.I3(CLBLM_R_X41Y100_SLICE_X67Y100_BQ),
.I4(CLBLL_L_X42Y107_SLICE_X69Y107_A5Q),
.I5(CLBLL_L_X42Y107_SLICE_X68Y107_BO5),
.O5(CLBLL_L_X42Y107_SLICE_X68Y107_AO5),
.O6(CLBLL_L_X42Y107_SLICE_X68Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y107_SLICE_X69Y107_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y107_SLICE_X69Y107_AO5),
.Q(CLBLL_L_X42Y107_SLICE_X69Y107_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y107_SLICE_X69Y107_B5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y107_SLICE_X69Y107_BO5),
.Q(CLBLL_L_X42Y107_SLICE_X69Y107_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y107_SLICE_X69Y107_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y107_SLICE_X69Y107_CO5),
.Q(CLBLL_L_X42Y107_SLICE_X69Y107_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y107_SLICE_X69Y107_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y107_SLICE_X69Y107_DO5),
.Q(CLBLL_L_X42Y107_SLICE_X69Y107_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y107_SLICE_X69Y107_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y112_SLICE_X68Y112_C5Q),
.Q(CLBLL_L_X42Y107_SLICE_X69Y107_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y107_SLICE_X69Y107_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y112_SLICE_X68Y112_CQ),
.Q(CLBLL_L_X42Y107_SLICE_X69Y107_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y107_SLICE_X69Y107_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y92_SLICE_X68Y92_BQ),
.Q(CLBLL_L_X42Y107_SLICE_X69Y107_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y107_SLICE_X69Y107_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y112_SLICE_X68Y112_A5Q),
.Q(CLBLL_L_X42Y107_SLICE_X69Y107_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaaaaaa)
  ) CLBLL_L_X42Y107_SLICE_X69Y107_DLUT (
.I0(CLBLL_L_X42Y112_SLICE_X68Y112_AQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y107_SLICE_X69Y107_DO5),
.O6(CLBLL_L_X42Y107_SLICE_X69Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLL_L_X42Y107_SLICE_X69Y107_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X42Y92_SLICE_X68Y92_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y107_SLICE_X69Y107_CO5),
.O6(CLBLL_L_X42Y107_SLICE_X69Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f0f0f0f0)
  ) CLBLL_L_X42Y107_SLICE_X69Y107_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y92_SLICE_X68Y92_D5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y107_SLICE_X69Y107_BO5),
.O6(CLBLL_L_X42Y107_SLICE_X69Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff0000)
  ) CLBLL_L_X42Y107_SLICE_X69Y107_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X42Y112_SLICE_X68Y112_B5Q),
.I5(1'b1),
.O5(CLBLL_L_X42Y107_SLICE_X69Y107_AO5),
.O6(CLBLL_L_X42Y107_SLICE_X69Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y108_SLICE_X68Y108_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y102_SLICE_X66Y102_AO5),
.D(CLBLL_L_X42Y108_SLICE_X68Y108_CO5),
.Q(CLBLL_L_X42Y108_SLICE_X68Y108_C5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fa72f0f0)
  ) CLBLL_L_X42Y108_SLICE_X68Y108_DLUT (
.I0(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I1(CLBLL_L_X42Y108_SLICE_X68Y108_C5Q),
.I2(CLBLL_L_X42Y68_SLICE_X68Y68_B5Q),
.I3(CLBLL_L_X42Y111_SLICE_X69Y111_A5Q),
.I4(CLBLL_L_X42Y109_SLICE_X69Y109_BO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y108_SLICE_X68Y108_DO5),
.O6(CLBLL_L_X42Y108_SLICE_X68Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000050505050)
  ) CLBLL_L_X42Y108_SLICE_X68Y108_CLUT (
.I0(CLBLL_L_X42Y102_SLICE_X68Y102_AO6),
.I1(1'b1),
.I2(CLBLL_L_X42Y109_SLICE_X69Y109_CO6),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y108_SLICE_X68Y108_CO5),
.O6(CLBLL_L_X42Y108_SLICE_X68Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000035551555)
  ) CLBLL_L_X42Y108_SLICE_X68Y108_BLUT (
.I0(CLBLL_L_X42Y105_SLICE_X69Y105_AQ),
.I1(CLBLL_L_X42Y111_SLICE_X69Y111_AQ),
.I2(CLBLL_L_X42Y109_SLICE_X69Y109_BO6),
.I3(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I4(CLBLL_L_X42Y108_SLICE_X68Y108_C5Q),
.I5(1'b1),
.O5(CLBLL_L_X42Y108_SLICE_X68Y108_BO5),
.O6(CLBLL_L_X42Y108_SLICE_X68Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fcf074f0)
  ) CLBLL_L_X42Y108_SLICE_X68Y108_ALUT (
.I0(CLBLL_L_X42Y108_SLICE_X68Y108_C5Q),
.I1(CLBLL_L_X42Y109_SLICE_X69Y109_BO6),
.I2(CLBLL_L_X42Y68_SLICE_X68Y68_D5Q),
.I3(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I4(CLBLL_L_X42Y111_SLICE_X69Y111_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y108_SLICE_X68Y108_AO5),
.O6(CLBLL_L_X42Y108_SLICE_X68Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y108_SLICE_X69Y108_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y108_SLICE_X69Y108_AO5),
.Q(CLBLL_L_X42Y108_SLICE_X69Y108_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y108_SLICE_X69Y108_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y108_SLICE_X69Y108_DO5),
.Q(CLBLL_L_X42Y108_SLICE_X69Y108_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y108_SLICE_X69Y108_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y111_SLICE_X68Y111_D5Q),
.Q(CLBLL_L_X42Y108_SLICE_X69Y108_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y108_SLICE_X69Y108_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y101_SLICE_X69Y101_CQ),
.Q(CLBLL_L_X42Y108_SLICE_X69Y108_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaaaaaa)
  ) CLBLL_L_X42Y108_SLICE_X69Y108_DLUT (
.I0(CLBLL_L_X42Y111_SLICE_X68Y111_C5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y108_SLICE_X69Y108_DO5),
.O6(CLBLL_L_X42Y108_SLICE_X69Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000fffe00fe)
  ) CLBLL_L_X42Y108_SLICE_X69Y108_CLUT (
.I0(CLBLM_R_X41Y102_SLICE_X66Y102_AO6),
.I1(CLBLM_R_X41Y108_SLICE_X67Y108_BO6),
.I2(CLBLL_L_X42Y102_SLICE_X68Y102_AO5),
.I3(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.I4(CLBLL_L_X42Y110_SLICE_X68Y110_BO5),
.I5(1'b1),
.O5(CLBLL_L_X42Y108_SLICE_X69Y108_CO5),
.O6(CLBLL_L_X42Y108_SLICE_X69Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000dc8ccccc)
  ) CLBLL_L_X42Y108_SLICE_X69Y108_BLUT (
.I0(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I1(CLBLL_L_X42Y108_SLICE_X69Y108_DQ),
.I2(CLBLM_R_X41Y108_SLICE_X67Y108_BO6),
.I3(CLBLL_L_X42Y108_SLICE_X69Y108_A5Q),
.I4(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y108_SLICE_X69Y108_BO5),
.O6(CLBLL_L_X42Y108_SLICE_X69Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLL_L_X42Y108_SLICE_X69Y108_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y111_SLICE_X68Y111_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y108_SLICE_X69Y108_AO5),
.O6(CLBLL_L_X42Y108_SLICE_X69Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y109_SLICE_X68Y109_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLL_L_X42Y109_SLICE_X68Y109_DO5),
.Q(CLBLL_L_X42Y109_SLICE_X68Y109_D5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y109_SLICE_X68Y109_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLM_R_X41Y108_SLICE_X66Y108_AO6),
.Q(CLBLL_L_X42Y109_SLICE_X68Y109_DQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0fcccccccc)
  ) CLBLL_L_X42Y109_SLICE_X68Y109_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y109_SLICE_X68Y109_AO6),
.I2(CLBLM_R_X41Y109_SLICE_X66Y109_BO5),
.I3(1'b1),
.I4(CLBLM_R_X41Y102_SLICE_X66Y102_AO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y109_SLICE_X68Y109_DO5),
.O6(CLBLL_L_X42Y109_SLICE_X68Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001000000000)
  ) CLBLL_L_X42Y109_SLICE_X68Y109_CLUT (
.I0(CLBLL_L_X42Y109_SLICE_X68Y109_D5Q),
.I1(CLBLM_R_X41Y108_SLICE_X66Y108_D5Q),
.I2(CLBLM_R_X41Y110_SLICE_X66Y110_AO6),
.I3(CLBLL_L_X42Y102_SLICE_X68Y102_BQ),
.I4(CLBLL_L_X42Y109_SLICE_X68Y109_DQ),
.I5(CLBLM_R_X41Y108_SLICE_X67Y108_CO5),
.O5(CLBLL_L_X42Y109_SLICE_X68Y109_CO5),
.O6(CLBLL_L_X42Y109_SLICE_X68Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000100000000)
  ) CLBLL_L_X42Y109_SLICE_X68Y109_BLUT (
.I0(CLBLM_R_X41Y102_SLICE_X67Y102_C5Q),
.I1(CLBLL_L_X42Y108_SLICE_X68Y108_C5Q),
.I2(CLBLL_L_X42Y109_SLICE_X69Y109_DQ),
.I3(CLBLL_L_X42Y102_SLICE_X68Y102_BQ),
.I4(CLBLL_L_X42Y109_SLICE_X68Y109_D5Q),
.I5(CLBLM_R_X41Y110_SLICE_X66Y110_AO6),
.O5(CLBLL_L_X42Y109_SLICE_X68Y109_BO5),
.O6(CLBLL_L_X42Y109_SLICE_X68Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000cffb30080)
  ) CLBLL_L_X42Y109_SLICE_X68Y109_ALUT (
.I0(CLBLL_L_X42Y110_SLICE_X69Y110_BO5),
.I1(CLBLL_L_X42Y109_SLICE_X68Y109_DO6),
.I2(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I3(CLBLM_R_X41Y115_SLICE_X66Y115_DO6),
.I4(CLBLL_L_X42Y109_SLICE_X68Y109_D5Q),
.I5(CLBLM_R_X41Y109_SLICE_X66Y109_CO6),
.O5(CLBLL_L_X42Y109_SLICE_X68Y109_AO5),
.O6(CLBLL_L_X42Y109_SLICE_X68Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y109_SLICE_X69Y109_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y110_SLICE_X69Y110_AO5),
.D(CLBLL_L_X42Y109_SLICE_X69Y109_DO6),
.Q(CLBLL_L_X42Y109_SLICE_X69Y109_DQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hccceccce00000000)
  ) CLBLL_L_X42Y109_SLICE_X69Y109_DLUT (
.I0(CLBLL_L_X42Y109_SLICE_X69Y109_DQ),
.I1(CLBLL_L_X42Y110_SLICE_X68Y110_AO5),
.I2(CLBLM_R_X41Y102_SLICE_X66Y102_CO6),
.I3(CLBLL_L_X42Y103_SLICE_X68Y103_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y109_SLICE_X69Y109_DO5),
.O6(CLBLL_L_X42Y109_SLICE_X69Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000c0055515115)
  ) CLBLL_L_X42Y109_SLICE_X69Y109_CLUT (
.I0(CLBLM_R_X41Y109_SLICE_X67Y109_CO6),
.I1(CLBLL_L_X42Y109_SLICE_X68Y109_CO6),
.I2(CLBLL_L_X42Y108_SLICE_X68Y108_C5Q),
.I3(CLBLM_R_X41Y102_SLICE_X67Y102_C5Q),
.I4(CLBLL_L_X42Y109_SLICE_X69Y109_DQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y109_SLICE_X69Y109_CO5),
.O6(CLBLL_L_X42Y109_SLICE_X69Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0303030300005500)
  ) CLBLL_L_X42Y109_SLICE_X69Y109_BLUT (
.I0(CLBLL_L_X42Y110_SLICE_X68Y110_AO5),
.I1(CLBLL_L_X42Y109_SLICE_X69Y109_DQ),
.I2(CLBLM_R_X41Y102_SLICE_X67Y102_C5Q),
.I3(CLBLL_L_X42Y109_SLICE_X69Y109_CO5),
.I4(CLBLM_R_X41Y109_SLICE_X67Y109_CO5),
.I5(1'b1),
.O5(CLBLL_L_X42Y109_SLICE_X69Y109_BO5),
.O6(CLBLL_L_X42Y109_SLICE_X69Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7070407070707070)
  ) CLBLL_L_X42Y109_SLICE_X69Y109_ALUT (
.I0(CLBLL_L_X42Y110_SLICE_X69Y110_AQ),
.I1(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(CLBLL_L_X42Y109_SLICE_X69Y109_BO5),
.I4(CLBLM_R_X41Y109_SLICE_X66Y109_CO6),
.I5(CLBLL_L_X42Y110_SLICE_X68Y110_DO5),
.O5(CLBLL_L_X42Y109_SLICE_X69Y109_AO5),
.O6(CLBLL_L_X42Y109_SLICE_X69Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y110_SLICE_X68Y110_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y110_SLICE_X68Y110_BO6),
.D(CLBLL_L_X42Y110_SLICE_X68Y110_CO5),
.Q(CLBLL_L_X42Y110_SLICE_X68Y110_C5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000333300f000f0)
  ) CLBLL_L_X42Y110_SLICE_X68Y110_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X41Y109_SLICE_X67Y109_BO6),
.I2(CLBLL_L_X42Y110_SLICE_X68Y110_DO6),
.I3(CLBLM_R_X41Y109_SLICE_X67Y109_BO5),
.I4(CLBLL_L_X42Y110_SLICE_X68Y110_AO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y110_SLICE_X68Y110_DO5),
.O6(CLBLL_L_X42Y110_SLICE_X68Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff8f0f)
  ) CLBLL_L_X42Y110_SLICE_X68Y110_CLUT (
.I0(CLBLL_L_X42Y110_SLICE_X68Y110_C5Q),
.I1(CLBLL_L_X42Y109_SLICE_X69Y109_BO5),
.I2(CLBLM_R_X41Y116_SLICE_X67Y116_BO5),
.I3(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I4(CLBLL_L_X42Y104_SLICE_X68Y104_BO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y110_SLICE_X68Y110_CO5),
.O6(CLBLL_L_X42Y110_SLICE_X68Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hff330f3388888888)
  ) CLBLL_L_X42Y110_SLICE_X68Y110_BLUT (
.I0(CLBLL_L_X42Y109_SLICE_X69Y109_CO5),
.I1(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I2(CLBLL_L_X42Y110_SLICE_X68Y110_DO5),
.I3(CLBLL_L_X42Y109_SLICE_X69Y109_BO5),
.I4(CLBLM_R_X41Y109_SLICE_X66Y109_CO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y110_SLICE_X68Y110_BO5),
.O6(CLBLL_L_X42Y110_SLICE_X68Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0080008020002000)
  ) CLBLL_L_X42Y110_SLICE_X68Y110_ALUT (
.I0(CLBLM_R_X41Y110_SLICE_X66Y110_AO6),
.I1(CLBLL_L_X42Y102_SLICE_X68Y102_BQ),
.I2(CLBLM_R_X41Y109_SLICE_X66Y109_DO5),
.I3(CLBLL_L_X42Y109_SLICE_X68Y109_D5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y110_SLICE_X68Y110_AO5),
.O6(CLBLL_L_X42Y110_SLICE_X68Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y110_SLICE_X69Y110_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLL_L_X42Y110_SLICE_X69Y110_CO5),
.Q(CLBLL_L_X42Y110_SLICE_X69Y110_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y110_SLICE_X69Y110_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLL_L_X42Y110_SLICE_X69Y110_DO5),
.Q(CLBLL_L_X42Y110_SLICE_X69Y110_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y110_SLICE_X69Y110_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLL_L_X42Y109_SLICE_X69Y109_AO6),
.Q(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000088808080)
  ) CLBLL_L_X42Y110_SLICE_X69Y110_DLUT (
.I0(CLBLL_L_X42Y71_SLICE_X68Y71_BQ),
.I1(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I2(CLBLL_L_X42Y110_SLICE_X69Y110_AQ),
.I3(CLBLL_L_X42Y112_SLICE_X69Y112_BQ),
.I4(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y110_SLICE_X69Y110_DO5),
.O6(CLBLL_L_X42Y110_SLICE_X69Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555662aaaaa)
  ) CLBLL_L_X42Y110_SLICE_X69Y110_CLUT (
.I0(CLBLL_L_X42Y110_SLICE_X69Y110_C5Q),
.I1(CLBLL_L_X42Y71_SLICE_X68Y71_BQ),
.I2(CLBLL_L_X42Y112_SLICE_X69Y112_DQ),
.I3(CLBLL_L_X42Y112_SLICE_X69Y112_C5Q),
.I4(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y110_SLICE_X69Y110_CO5),
.O6(CLBLL_L_X42Y110_SLICE_X69Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0088000022000000)
  ) CLBLL_L_X42Y110_SLICE_X69Y110_BLUT (
.I0(CLBLM_R_X41Y109_SLICE_X66Y109_DO5),
.I1(CLBLL_L_X42Y102_SLICE_X68Y102_BQ),
.I2(1'b1),
.I3(CLBLL_L_X42Y109_SLICE_X68Y109_D5Q),
.I4(CLBLM_R_X41Y110_SLICE_X66Y110_AO6),
.I5(1'b1),
.O5(CLBLL_L_X42Y110_SLICE_X69Y110_BO5),
.O6(CLBLL_L_X42Y110_SLICE_X69Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000002220222)
  ) CLBLL_L_X42Y110_SLICE_X69Y110_ALUT (
.I0(CLBLL_L_X42Y109_SLICE_X68Y109_DO6),
.I1(CLBLM_R_X41Y115_SLICE_X66Y115_DO6),
.I2(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I3(CLBLL_L_X42Y110_SLICE_X69Y110_BO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y110_SLICE_X69Y110_AO5),
.O6(CLBLL_L_X42Y110_SLICE_X69Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y111_SLICE_X68Y111_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(BRAM_L_X44Y95_RAMB18_X2Y38_DO7),
.Q(CLBLL_L_X42Y111_SLICE_X68Y111_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y111_SLICE_X68Y111_B5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(BRAM_L_X44Y95_RAMB18_X2Y38_DO2),
.Q(CLBLL_L_X42Y111_SLICE_X68Y111_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y111_SLICE_X68Y111_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(BRAM_L_X44Y95_RAMB18_X2Y38_DO4),
.Q(CLBLL_L_X42Y111_SLICE_X68Y111_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y111_SLICE_X68Y111_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y94_SLICE_X68Y94_BQ),
.Q(CLBLL_L_X42Y111_SLICE_X68Y111_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y111_SLICE_X68Y111_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y111_SLICE_X68Y111_AO5),
.Q(CLBLL_L_X42Y111_SLICE_X68Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y111_SLICE_X68Y111_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y111_SLICE_X68Y111_BO5),
.Q(CLBLL_L_X42Y111_SLICE_X68Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y111_SLICE_X68Y111_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y111_SLICE_X68Y111_CO5),
.Q(CLBLL_L_X42Y111_SLICE_X68Y111_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y111_SLICE_X68Y111_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y111_SLICE_X68Y111_DO5),
.Q(CLBLL_L_X42Y111_SLICE_X68Y111_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLL_L_X42Y111_SLICE_X68Y111_DLUT (
.I0(1'b1),
.I1(BRAM_L_X44Y95_RAMB18_X2Y38_DO5),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y111_SLICE_X68Y111_DO5),
.O6(CLBLL_L_X42Y111_SLICE_X68Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLL_L_X42Y111_SLICE_X68Y111_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_L_X44Y95_RAMB18_X2Y38_DO10),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y111_SLICE_X68Y111_CO5),
.O6(CLBLL_L_X42Y111_SLICE_X68Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff0000)
  ) CLBLL_L_X42Y111_SLICE_X68Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(BRAM_L_X44Y95_RAMB18_X2Y38_DOP0),
.I5(1'b1),
.O5(CLBLL_L_X42Y111_SLICE_X68Y111_BO5),
.O6(CLBLL_L_X42Y111_SLICE_X68Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLL_L_X42Y111_SLICE_X68Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(BRAM_L_X44Y95_RAMB18_X2Y38_DO9),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y111_SLICE_X68Y111_AO5),
.O6(CLBLL_L_X42Y111_SLICE_X68Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y111_SLICE_X69Y111_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y111_SLICE_X69Y111_AO5),
.Q(CLBLL_L_X42Y111_SLICE_X69Y111_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y111_SLICE_X69Y111_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y111_SLICE_X69Y111_DO5),
.Q(CLBLL_L_X42Y111_SLICE_X69Y111_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y111_SLICE_X69Y111_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y111_SLICE_X68Y111_A5Q),
.Q(CLBLL_L_X42Y111_SLICE_X69Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y111_SLICE_X69Y111_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y98_SLICE_X69Y98_BQ),
.Q(CLBLL_L_X42Y111_SLICE_X69Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y111_SLICE_X69Y111_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y111_SLICE_X68Y111_AQ),
.Q(CLBLL_L_X42Y111_SLICE_X69Y111_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLL_L_X42Y111_SLICE_X69Y111_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y111_SLICE_X68Y111_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y111_SLICE_X69Y111_DO5),
.O6(CLBLL_L_X42Y111_SLICE_X69Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000f0f5511)
  ) CLBLL_L_X42Y111_SLICE_X69Y111_CLUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_DO6),
.I1(CLBLM_R_X41Y106_SLICE_X67Y106_BO5),
.I2(CLBLL_L_X42Y105_SLICE_X69Y105_BO5),
.I3(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I4(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y111_SLICE_X69Y111_CO5),
.O6(CLBLL_L_X42Y111_SLICE_X69Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y111_SLICE_X69Y111_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y111_SLICE_X69Y111_BO5),
.O6(CLBLL_L_X42Y111_SLICE_X69Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLL_L_X42Y111_SLICE_X69Y111_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y111_SLICE_X68Y111_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y111_SLICE_X69Y111_AO5),
.O6(CLBLL_L_X42Y111_SLICE_X69Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y112_SLICE_X68Y112_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y91_SLICE_X68Y91_AQ),
.Q(CLBLL_L_X42Y112_SLICE_X68Y112_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y112_SLICE_X68Y112_B5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y90_SLICE_X68Y90_AQ),
.Q(CLBLL_L_X42Y112_SLICE_X68Y112_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y112_SLICE_X68Y112_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y90_SLICE_X68Y90_BQ),
.Q(CLBLL_L_X42Y112_SLICE_X68Y112_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y112_SLICE_X68Y112_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y113_SLICE_X68Y113_D5Q),
.Q(CLBLL_L_X42Y112_SLICE_X68Y112_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y112_SLICE_X68Y112_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y112_SLICE_X68Y112_AO5),
.Q(CLBLL_L_X42Y112_SLICE_X68Y112_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y112_SLICE_X68Y112_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y112_SLICE_X68Y112_BO5),
.Q(CLBLL_L_X42Y112_SLICE_X68Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y112_SLICE_X68Y112_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y112_SLICE_X68Y112_CO5),
.Q(CLBLL_L_X42Y112_SLICE_X68Y112_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y112_SLICE_X68Y112_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y112_SLICE_X68Y112_DO5),
.Q(CLBLL_L_X42Y112_SLICE_X68Y112_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLL_L_X42Y112_SLICE_X68Y112_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y90_SLICE_X68Y90_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y112_SLICE_X68Y112_DO5),
.O6(CLBLL_L_X42Y112_SLICE_X68Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLL_L_X42Y112_SLICE_X68Y112_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X42Y91_SLICE_X68Y91_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y112_SLICE_X68Y112_CO5),
.O6(CLBLL_L_X42Y112_SLICE_X68Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff0000)
  ) CLBLL_L_X42Y112_SLICE_X68Y112_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X42Y91_SLICE_X68Y91_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y112_SLICE_X68Y112_BO5),
.O6(CLBLL_L_X42Y112_SLICE_X68Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLL_L_X42Y112_SLICE_X68Y112_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X42Y91_SLICE_X68Y91_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y112_SLICE_X68Y112_AO5),
.O6(CLBLL_L_X42Y112_SLICE_X68Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y112_SLICE_X69Y112_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLL_L_X42Y112_SLICE_X69Y112_CO5),
.Q(CLBLL_L_X42Y112_SLICE_X69Y112_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y112_SLICE_X69Y112_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLL_L_X42Y112_SLICE_X69Y112_AO6),
.Q(CLBLL_L_X42Y112_SLICE_X69Y112_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y112_SLICE_X69Y112_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLL_L_X42Y112_SLICE_X69Y112_BO5),
.Q(CLBLL_L_X42Y112_SLICE_X69Y112_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000080800000)
  ) CLBLL_L_X42Y112_SLICE_X69Y112_DLUT (
.I0(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I1(CLBLL_L_X42Y112_SLICE_X69Y112_BQ),
.I2(CLBLL_L_X42Y71_SLICE_X68Y71_BQ),
.I3(1'b1),
.I4(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y112_SLICE_X69Y112_DO5),
.O6(CLBLL_L_X42Y112_SLICE_X69Y112_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000c4c0cc00)
  ) CLBLL_L_X42Y112_SLICE_X69Y112_CLUT (
.I0(CLBLL_L_X42Y43_SLICE_X68Y43_D_XOR),
.I1(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I2(CLBLL_L_X42Y112_SLICE_X69Y112_DQ),
.I3(CLBLL_L_X42Y112_SLICE_X69Y112_C5Q),
.I4(CLBLL_L_X42Y71_SLICE_X68Y71_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y112_SLICE_X69Y112_CO5),
.O6(CLBLL_L_X42Y112_SLICE_X69Y112_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff88)
  ) CLBLL_L_X42Y112_SLICE_X69Y112_BLUT (
.I0(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I1(CLBLL_L_X42Y112_SLICE_X69Y112_DQ),
.I2(1'b1),
.I3(CLBLL_L_X42Y112_SLICE_X69Y112_DO5),
.I4(CLBLL_L_X42Y71_SLICE_X68Y71_BQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y112_SLICE_X69Y112_BO5),
.O6(CLBLL_L_X42Y112_SLICE_X69Y112_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfdfd75f575f575f5)
  ) CLBLL_L_X42Y112_SLICE_X69Y112_ALUT (
.I0(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I1(CLBLL_L_X42Y71_SLICE_X68Y71_BQ),
.I2(CLBLL_L_X42Y112_SLICE_X69Y112_BQ),
.I3(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I4(CLBLL_L_X42Y112_SLICE_X69Y112_C5Q),
.I5(CLBLL_L_X42Y43_SLICE_X68Y43_D_XOR),
.O5(CLBLL_L_X42Y112_SLICE_X69Y112_AO5),
.O6(CLBLL_L_X42Y112_SLICE_X69Y112_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y113_SLICE_X68Y113_D5_FDSE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y96_SLICE_X68Y96_CO5),
.D(CLBLL_L_X42Y96_SLICE_X68Y96_BO6),
.Q(CLBLL_L_X42Y113_SLICE_X68Y113_D5Q),
.S(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y113_SLICE_X68Y113_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y113_SLICE_X68Y113_DO5),
.O6(CLBLL_L_X42Y113_SLICE_X68Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y113_SLICE_X68Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y113_SLICE_X68Y113_CO5),
.O6(CLBLL_L_X42Y113_SLICE_X68Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y113_SLICE_X68Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y113_SLICE_X68Y113_BO5),
.O6(CLBLL_L_X42Y113_SLICE_X68Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y113_SLICE_X68Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y113_SLICE_X68Y113_AO5),
.O6(CLBLL_L_X42Y113_SLICE_X68Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y113_SLICE_X69Y113_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y93_SLICE_X68Y93_BQ),
.Q(CLBLL_L_X42Y113_SLICE_X69Y113_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y113_SLICE_X69Y113_B5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y97_SLICE_X68Y97_AQ),
.Q(CLBLL_L_X42Y113_SLICE_X69Y113_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y113_SLICE_X69Y113_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y104_SLICE_X69Y104_CQ),
.Q(CLBLL_L_X42Y113_SLICE_X69Y113_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y113_SLICE_X69Y113_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y104_SLICE_X69Y104_BQ),
.Q(CLBLL_L_X42Y113_SLICE_X69Y113_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y113_SLICE_X69Y113_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y113_SLICE_X69Y113_AO5),
.Q(CLBLL_L_X42Y113_SLICE_X69Y113_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y113_SLICE_X69Y113_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y113_SLICE_X69Y113_BO5),
.Q(CLBLL_L_X42Y113_SLICE_X69Y113_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y113_SLICE_X69Y113_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y113_SLICE_X69Y113_CO5),
.Q(CLBLL_L_X42Y113_SLICE_X69Y113_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y113_SLICE_X69Y113_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y97_SLICE_X69Y97_CO6),
.D(CLBLL_L_X42Y113_SLICE_X69Y113_DO5),
.Q(CLBLL_L_X42Y113_SLICE_X69Y113_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLL_L_X42Y113_SLICE_X69Y113_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y104_SLICE_X69Y104_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y113_SLICE_X69Y113_DO5),
.O6(CLBLL_L_X42Y113_SLICE_X69Y113_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLL_L_X42Y113_SLICE_X69Y113_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X42Y93_SLICE_X69Y93_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y113_SLICE_X69Y113_CO5),
.O6(CLBLL_L_X42Y113_SLICE_X69Y113_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff0000)
  ) CLBLL_L_X42Y113_SLICE_X69Y113_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X42Y93_SLICE_X68Y93_DQ),
.I5(1'b1),
.O5(CLBLL_L_X42Y113_SLICE_X69Y113_BO5),
.O6(CLBLL_L_X42Y113_SLICE_X69Y113_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLL_L_X42Y113_SLICE_X69Y113_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLL_L_X42Y93_SLICE_X68Y93_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y113_SLICE_X69Y113_AO5),
.O6(CLBLL_L_X42Y113_SLICE_X69Y113_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y118_SLICE_X68Y118_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y118_SLICE_X68Y118_DO5),
.O6(CLBLL_L_X42Y118_SLICE_X68Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y118_SLICE_X68Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y118_SLICE_X68Y118_CO5),
.O6(CLBLL_L_X42Y118_SLICE_X68Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y118_SLICE_X68Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y118_SLICE_X68Y118_BO5),
.O6(CLBLL_L_X42Y118_SLICE_X68Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X42Y118_SLICE_X68Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y118_SLICE_X68Y118_AO5),
.O6(CLBLL_L_X42Y118_SLICE_X68Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y118_SLICE_X69Y118_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y112_SLICE_X69Y112_DO5),
.D(CLBLL_L_X42Y118_SLICE_X69Y118_AO5),
.Q(CLBLL_L_X42Y118_SLICE_X69Y118_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y118_SLICE_X69Y118_B5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y112_SLICE_X69Y112_DO5),
.D(CLBLL_L_X42Y118_SLICE_X69Y118_BO5),
.Q(CLBLL_L_X42Y118_SLICE_X69Y118_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y118_SLICE_X69Y118_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y112_SLICE_X69Y112_DO5),
.D(CLBLL_L_X42Y118_SLICE_X69Y118_CO5),
.Q(CLBLL_L_X42Y118_SLICE_X69Y118_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y118_SLICE_X69Y118_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y112_SLICE_X69Y112_DO5),
.D(CLBLL_L_X42Y118_SLICE_X69Y118_DO5),
.Q(CLBLL_L_X42Y118_SLICE_X69Y118_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y118_SLICE_X69Y118_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y112_SLICE_X69Y112_DO5),
.D(CLBLM_R_X41Y105_SLICE_X66Y105_DQ),
.Q(CLBLL_L_X42Y118_SLICE_X69Y118_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y118_SLICE_X69Y118_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y112_SLICE_X69Y112_DO5),
.D(CLBLM_R_X41Y103_SLICE_X67Y103_D5Q),
.Q(CLBLL_L_X42Y118_SLICE_X69Y118_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y118_SLICE_X69Y118_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y112_SLICE_X69Y112_DO5),
.D(CLBLM_R_X41Y104_SLICE_X67Y104_C5Q),
.Q(CLBLL_L_X42Y118_SLICE_X69Y118_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X42Y118_SLICE_X69Y118_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y112_SLICE_X69Y112_DO5),
.D(CLBLM_R_X41Y110_SLICE_X67Y110_B5Q),
.Q(CLBLL_L_X42Y118_SLICE_X69Y118_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaaaaaa)
  ) CLBLL_L_X42Y118_SLICE_X69Y118_DLUT (
.I0(CLBLL_L_X42Y110_SLICE_X68Y110_C5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y118_SLICE_X69Y118_DO5),
.O6(CLBLL_L_X42Y118_SLICE_X69Y118_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLL_L_X42Y118_SLICE_X69Y118_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X41Y107_SLICE_X67Y107_D5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y118_SLICE_X69Y118_CO5),
.O6(CLBLL_L_X42Y118_SLICE_X69Y118_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f0f0f0f0)
  ) CLBLL_L_X42Y118_SLICE_X69Y118_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X41Y104_SLICE_X66Y104_D5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X42Y118_SLICE_X69Y118_BO5),
.O6(CLBLL_L_X42Y118_SLICE_X69Y118_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff0000)
  ) CLBLL_L_X42Y118_SLICE_X69Y118_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X41Y111_SLICE_X67Y111_A5Q),
.I5(1'b1),
.O5(CLBLL_L_X42Y118_SLICE_X69Y118_AO5),
.O6(CLBLL_L_X42Y118_SLICE_X69Y118_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y54_SLICE_X2Y54_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y54_SLICE_X2Y54_DO5),
.O6(CLBLM_R_X3Y54_SLICE_X2Y54_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y54_SLICE_X2Y54_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y54_SLICE_X2Y54_CO5),
.O6(CLBLM_R_X3Y54_SLICE_X2Y54_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y54_SLICE_X2Y54_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y54_SLICE_X2Y54_BO5),
.O6(CLBLM_R_X3Y54_SLICE_X2Y54_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y54_SLICE_X2Y54_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y54_SLICE_X2Y54_AO5),
.O6(CLBLM_R_X3Y54_SLICE_X2Y54_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y54_SLICE_X3Y54_B5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y54_SLICE_X3Y54_BO5),
.Q(CLBLM_R_X3Y54_SLICE_X3Y54_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y54_SLICE_X3Y54_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y54_SLICE_X3Y54_B_XOR),
.Q(CLBLM_R_X3Y54_SLICE_X3Y54_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y54_SLICE_X3Y54_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y54_SLICE_X3Y54_C_XOR),
.Q(CLBLM_R_X3Y54_SLICE_X3Y54_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y54_SLICE_X3Y54_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y54_SLICE_X3Y54_D_XOR),
.Q(CLBLM_R_X3Y54_SLICE_X3Y54_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y54_SLICE_X3Y54_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X3Y54_SLICE_X3Y54_D_CY, CLBLM_R_X3Y54_SLICE_X3Y54_C_CY, CLBLM_R_X3Y54_SLICE_X3Y54_B_CY, CLBLM_R_X3Y54_SLICE_X3Y54_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({CLBLM_R_X3Y54_SLICE_X3Y54_D_XOR, CLBLM_R_X3Y54_SLICE_X3Y54_C_XOR, CLBLM_R_X3Y54_SLICE_X3Y54_B_XOR, CLBLM_R_X3Y54_SLICE_X3Y54_A_XOR}),
.S({CLBLM_R_X3Y54_SLICE_X3Y54_DO6, CLBLM_R_X3Y54_SLICE_X3Y54_CO6, CLBLM_R_X3Y54_SLICE_X3Y54_BO6, CLBLM_R_X3Y54_SLICE_X3Y54_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000000000)
  ) CLBLM_R_X3Y54_SLICE_X3Y54_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y54_SLICE_X3Y54_DQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y54_SLICE_X3Y54_DO5),
.O6(CLBLM_R_X3Y54_SLICE_X3Y54_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLM_R_X3Y54_SLICE_X3Y54_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y54_SLICE_X3Y54_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y54_SLICE_X3Y54_CO5),
.O6(CLBLM_R_X3Y54_SLICE_X3Y54_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000cccccccc)
  ) CLBLM_R_X3Y54_SLICE_X3Y54_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y54_SLICE_X3Y54_AO5),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y54_SLICE_X3Y54_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y54_SLICE_X3Y54_BO5),
.O6(CLBLM_R_X3Y54_SLICE_X3Y54_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000f0f0f0f)
  ) CLBLM_R_X3Y54_SLICE_X3Y54_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y54_SLICE_X3Y54_B5Q),
.I3(CLBLM_R_X3Y54_SLICE_X3Y54_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y54_SLICE_X3Y54_AO5),
.O6(CLBLM_R_X3Y54_SLICE_X3Y54_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y55_SLICE_X2Y55_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y55_SLICE_X2Y55_DO5),
.O6(CLBLM_R_X3Y55_SLICE_X2Y55_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y55_SLICE_X2Y55_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y55_SLICE_X2Y55_CO5),
.O6(CLBLM_R_X3Y55_SLICE_X2Y55_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y55_SLICE_X2Y55_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y55_SLICE_X2Y55_BO5),
.O6(CLBLM_R_X3Y55_SLICE_X2Y55_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y55_SLICE_X2Y55_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y55_SLICE_X2Y55_AO5),
.O6(CLBLM_R_X3Y55_SLICE_X2Y55_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y55_SLICE_X3Y55_B5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y55_SLICE_X3Y55_BO5),
.Q(CLBLM_R_X3Y55_SLICE_X3Y55_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y55_SLICE_X3Y55_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y55_SLICE_X3Y55_AO5),
.Q(CLBLM_R_X3Y55_SLICE_X3Y55_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y55_SLICE_X3Y55_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y55_SLICE_X3Y55_B_XOR),
.Q(CLBLM_R_X3Y55_SLICE_X3Y55_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y55_SLICE_X3Y55_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y55_SLICE_X3Y55_DO5),
.Q(CLBLM_R_X3Y55_SLICE_X3Y55_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y55_SLICE_X3Y55_CARRY4 (
.CI(CLBLM_R_X3Y54_SLICE_X3Y54_COUT),
.CO({CLBLM_R_X3Y55_SLICE_X3Y55_COUT, CLBLM_R_X3Y55_SLICE_X3Y55_C_CY, CLBLM_R_X3Y55_SLICE_X3Y55_B_CY, CLBLM_R_X3Y55_SLICE_X3Y55_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X3Y55_SLICE_X3Y55_D_XOR, CLBLM_R_X3Y55_SLICE_X3Y55_C_XOR, CLBLM_R_X3Y55_SLICE_X3Y55_B_XOR, CLBLM_R_X3Y55_SLICE_X3Y55_A_XOR}),
.S({CLBLM_R_X3Y55_SLICE_X3Y55_DO6, CLBLM_R_X3Y55_SLICE_X3Y55_CO6, CLBLM_R_X3Y55_SLICE_X3Y55_BO6, CLBLM_R_X3Y55_SLICE_X3Y55_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X3Y55_SLICE_X3Y55_DLUT (
.I0(CLBLM_R_X3Y55_SLICE_X3Y55_C_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y55_SLICE_X3Y55_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y55_SLICE_X3Y55_DO5),
.O6(CLBLM_R_X3Y55_SLICE_X3Y55_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLM_R_X3Y55_SLICE_X3Y55_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y55_SLICE_X3Y55_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y55_SLICE_X3Y55_CO5),
.O6(CLBLM_R_X3Y55_SLICE_X3Y55_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLM_R_X3Y55_SLICE_X3Y55_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y55_SLICE_X3Y55_BQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y55_SLICE_X3Y55_A_XOR),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y55_SLICE_X3Y55_BO5),
.O6(CLBLM_R_X3Y55_SLICE_X3Y55_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X3Y55_SLICE_X3Y55_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y55_SLICE_X3Y55_B5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y55_SLICE_X3Y55_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X3Y55_SLICE_X3Y55_AO5),
.O6(CLBLM_R_X3Y55_SLICE_X3Y55_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y56_SLICE_X2Y56_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y56_SLICE_X2Y56_DO5),
.O6(CLBLM_R_X3Y56_SLICE_X2Y56_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y56_SLICE_X2Y56_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y56_SLICE_X2Y56_CO5),
.O6(CLBLM_R_X3Y56_SLICE_X2Y56_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y56_SLICE_X2Y56_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y56_SLICE_X2Y56_BO5),
.O6(CLBLM_R_X3Y56_SLICE_X2Y56_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y56_SLICE_X2Y56_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y56_SLICE_X2Y56_AO5),
.O6(CLBLM_R_X3Y56_SLICE_X2Y56_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y56_SLICE_X3Y56_B5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y56_SLICE_X3Y56_BO5),
.Q(CLBLM_R_X3Y56_SLICE_X3Y56_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y56_SLICE_X3Y56_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y56_SLICE_X3Y56_AO5),
.Q(CLBLM_R_X3Y56_SLICE_X3Y56_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y56_SLICE_X3Y56_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y56_SLICE_X3Y56_B_XOR),
.Q(CLBLM_R_X3Y56_SLICE_X3Y56_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y56_SLICE_X3Y56_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y56_SLICE_X3Y56_DO5),
.Q(CLBLM_R_X3Y56_SLICE_X3Y56_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y56_SLICE_X3Y56_CARRY4 (
.CI(CLBLM_R_X3Y55_SLICE_X3Y55_COUT),
.CO({CLBLM_R_X3Y56_SLICE_X3Y56_COUT, CLBLM_R_X3Y56_SLICE_X3Y56_C_CY, CLBLM_R_X3Y56_SLICE_X3Y56_B_CY, CLBLM_R_X3Y56_SLICE_X3Y56_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X3Y56_SLICE_X3Y56_D_XOR, CLBLM_R_X3Y56_SLICE_X3Y56_C_XOR, CLBLM_R_X3Y56_SLICE_X3Y56_B_XOR, CLBLM_R_X3Y56_SLICE_X3Y56_A_XOR}),
.S({CLBLM_R_X3Y56_SLICE_X3Y56_DO6, CLBLM_R_X3Y56_SLICE_X3Y56_CO6, CLBLM_R_X3Y56_SLICE_X3Y56_BO6, CLBLM_R_X3Y56_SLICE_X3Y56_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X3Y56_SLICE_X3Y56_DLUT (
.I0(CLBLM_R_X3Y56_SLICE_X3Y56_C_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y56_SLICE_X3Y56_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y56_SLICE_X3Y56_DO5),
.O6(CLBLM_R_X3Y56_SLICE_X3Y56_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLM_R_X3Y56_SLICE_X3Y56_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y56_SLICE_X3Y56_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y56_SLICE_X3Y56_CO5),
.O6(CLBLM_R_X3Y56_SLICE_X3Y56_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLM_R_X3Y56_SLICE_X3Y56_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y56_SLICE_X3Y56_BQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y56_SLICE_X3Y56_A_XOR),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y56_SLICE_X3Y56_BO5),
.O6(CLBLM_R_X3Y56_SLICE_X3Y56_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X3Y56_SLICE_X3Y56_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y56_SLICE_X3Y56_B5Q),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y56_SLICE_X3Y56_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X3Y56_SLICE_X3Y56_AO5),
.O6(CLBLM_R_X3Y56_SLICE_X3Y56_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y57_SLICE_X2Y57_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y57_SLICE_X2Y57_DO5),
.O6(CLBLM_R_X3Y57_SLICE_X2Y57_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y57_SLICE_X2Y57_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y57_SLICE_X2Y57_CO5),
.O6(CLBLM_R_X3Y57_SLICE_X2Y57_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y57_SLICE_X2Y57_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y57_SLICE_X2Y57_BO5),
.O6(CLBLM_R_X3Y57_SLICE_X2Y57_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y57_SLICE_X2Y57_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y57_SLICE_X2Y57_AO5),
.O6(CLBLM_R_X3Y57_SLICE_X2Y57_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y57_SLICE_X3Y57_B5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y57_SLICE_X3Y57_BO5),
.Q(CLBLM_R_X3Y57_SLICE_X3Y57_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y57_SLICE_X3Y57_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y57_SLICE_X3Y57_AO5),
.Q(CLBLM_R_X3Y57_SLICE_X3Y57_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y57_SLICE_X3Y57_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y57_SLICE_X3Y57_B_XOR),
.Q(CLBLM_R_X3Y57_SLICE_X3Y57_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y57_SLICE_X3Y57_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y57_SLICE_X3Y57_DO5),
.Q(CLBLM_R_X3Y57_SLICE_X3Y57_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y57_SLICE_X3Y57_CARRY4 (
.CI(CLBLM_R_X3Y56_SLICE_X3Y56_COUT),
.CO({CLBLM_R_X3Y57_SLICE_X3Y57_COUT, CLBLM_R_X3Y57_SLICE_X3Y57_C_CY, CLBLM_R_X3Y57_SLICE_X3Y57_B_CY, CLBLM_R_X3Y57_SLICE_X3Y57_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X3Y57_SLICE_X3Y57_D_XOR, CLBLM_R_X3Y57_SLICE_X3Y57_C_XOR, CLBLM_R_X3Y57_SLICE_X3Y57_B_XOR, CLBLM_R_X3Y57_SLICE_X3Y57_A_XOR}),
.S({CLBLM_R_X3Y57_SLICE_X3Y57_DO6, CLBLM_R_X3Y57_SLICE_X3Y57_CO6, CLBLM_R_X3Y57_SLICE_X3Y57_BO6, CLBLM_R_X3Y57_SLICE_X3Y57_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X3Y57_SLICE_X3Y57_DLUT (
.I0(CLBLM_R_X3Y57_SLICE_X3Y57_A_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y57_SLICE_X3Y57_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y57_SLICE_X3Y57_DO5),
.O6(CLBLM_R_X3Y57_SLICE_X3Y57_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLM_R_X3Y57_SLICE_X3Y57_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y57_SLICE_X3Y57_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y57_SLICE_X3Y57_CO5),
.O6(CLBLM_R_X3Y57_SLICE_X3Y57_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X3Y57_SLICE_X3Y57_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y57_SLICE_X3Y57_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y57_SLICE_X3Y57_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X3Y57_SLICE_X3Y57_BO5),
.O6(CLBLM_R_X3Y57_SLICE_X3Y57_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X3Y57_SLICE_X3Y57_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y57_SLICE_X3Y57_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y57_SLICE_X3Y57_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X3Y57_SLICE_X3Y57_AO5),
.O6(CLBLM_R_X3Y57_SLICE_X3Y57_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y58_SLICE_X2Y58_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y58_SLICE_X2Y58_DO5),
.O6(CLBLM_R_X3Y58_SLICE_X2Y58_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y58_SLICE_X2Y58_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y58_SLICE_X2Y58_CO5),
.O6(CLBLM_R_X3Y58_SLICE_X2Y58_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y58_SLICE_X2Y58_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y58_SLICE_X2Y58_BO5),
.O6(CLBLM_R_X3Y58_SLICE_X2Y58_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y58_SLICE_X2Y58_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y58_SLICE_X2Y58_AO5),
.O6(CLBLM_R_X3Y58_SLICE_X2Y58_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y58_SLICE_X3Y58_B5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y58_SLICE_X3Y58_BO5),
.Q(CLBLM_R_X3Y58_SLICE_X3Y58_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y58_SLICE_X3Y58_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y58_SLICE_X3Y58_AO5),
.Q(CLBLM_R_X3Y58_SLICE_X3Y58_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y58_SLICE_X3Y58_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y58_SLICE_X3Y58_B_XOR),
.Q(CLBLM_R_X3Y58_SLICE_X3Y58_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y58_SLICE_X3Y58_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y58_SLICE_X3Y58_DO5),
.Q(CLBLM_R_X3Y58_SLICE_X3Y58_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y58_SLICE_X3Y58_CARRY4 (
.CI(CLBLM_R_X3Y57_SLICE_X3Y57_COUT),
.CO({CLBLM_R_X3Y58_SLICE_X3Y58_COUT, CLBLM_R_X3Y58_SLICE_X3Y58_C_CY, CLBLM_R_X3Y58_SLICE_X3Y58_B_CY, CLBLM_R_X3Y58_SLICE_X3Y58_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X3Y58_SLICE_X3Y58_D_XOR, CLBLM_R_X3Y58_SLICE_X3Y58_C_XOR, CLBLM_R_X3Y58_SLICE_X3Y58_B_XOR, CLBLM_R_X3Y58_SLICE_X3Y58_A_XOR}),
.S({CLBLM_R_X3Y58_SLICE_X3Y58_DO6, CLBLM_R_X3Y58_SLICE_X3Y58_CO6, CLBLM_R_X3Y58_SLICE_X3Y58_BO6, CLBLM_R_X3Y58_SLICE_X3Y58_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X3Y58_SLICE_X3Y58_DLUT (
.I0(CLBLM_R_X3Y58_SLICE_X3Y58_A_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y58_SLICE_X3Y58_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y58_SLICE_X3Y58_DO5),
.O6(CLBLM_R_X3Y58_SLICE_X3Y58_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLM_R_X3Y58_SLICE_X3Y58_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y58_SLICE_X3Y58_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y58_SLICE_X3Y58_CO5),
.O6(CLBLM_R_X3Y58_SLICE_X3Y58_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X3Y58_SLICE_X3Y58_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y58_SLICE_X3Y58_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y58_SLICE_X3Y58_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X3Y58_SLICE_X3Y58_BO5),
.O6(CLBLM_R_X3Y58_SLICE_X3Y58_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X3Y58_SLICE_X3Y58_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y58_SLICE_X3Y58_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y58_SLICE_X3Y58_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X3Y58_SLICE_X3Y58_AO5),
.O6(CLBLM_R_X3Y58_SLICE_X3Y58_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y59_SLICE_X2Y59_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y59_SLICE_X2Y59_DO5),
.O6(CLBLM_R_X3Y59_SLICE_X2Y59_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y59_SLICE_X2Y59_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y59_SLICE_X2Y59_CO5),
.O6(CLBLM_R_X3Y59_SLICE_X2Y59_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y59_SLICE_X2Y59_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y59_SLICE_X2Y59_BO5),
.O6(CLBLM_R_X3Y59_SLICE_X2Y59_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y59_SLICE_X2Y59_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y59_SLICE_X2Y59_AO5),
.O6(CLBLM_R_X3Y59_SLICE_X2Y59_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y59_SLICE_X3Y59_B5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y59_SLICE_X3Y59_BO5),
.Q(CLBLM_R_X3Y59_SLICE_X3Y59_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y59_SLICE_X3Y59_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y59_SLICE_X3Y59_AO5),
.Q(CLBLM_R_X3Y59_SLICE_X3Y59_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y59_SLICE_X3Y59_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y59_SLICE_X3Y59_B_XOR),
.Q(CLBLM_R_X3Y59_SLICE_X3Y59_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y59_SLICE_X3Y59_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y59_SLICE_X3Y59_DO5),
.Q(CLBLM_R_X3Y59_SLICE_X3Y59_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y59_SLICE_X3Y59_CARRY4 (
.CI(CLBLM_R_X3Y58_SLICE_X3Y58_COUT),
.CO({CLBLM_R_X3Y59_SLICE_X3Y59_COUT, CLBLM_R_X3Y59_SLICE_X3Y59_C_CY, CLBLM_R_X3Y59_SLICE_X3Y59_B_CY, CLBLM_R_X3Y59_SLICE_X3Y59_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X3Y59_SLICE_X3Y59_D_XOR, CLBLM_R_X3Y59_SLICE_X3Y59_C_XOR, CLBLM_R_X3Y59_SLICE_X3Y59_B_XOR, CLBLM_R_X3Y59_SLICE_X3Y59_A_XOR}),
.S({CLBLM_R_X3Y59_SLICE_X3Y59_DO6, CLBLM_R_X3Y59_SLICE_X3Y59_CO6, CLBLM_R_X3Y59_SLICE_X3Y59_BO6, CLBLM_R_X3Y59_SLICE_X3Y59_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ff00)
  ) CLBLM_R_X3Y59_SLICE_X3Y59_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y59_SLICE_X3Y59_B5Q),
.I3(CLBLM_R_X3Y59_SLICE_X3Y59_A_XOR),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y59_SLICE_X3Y59_DO5),
.O6(CLBLM_R_X3Y59_SLICE_X3Y59_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X3Y59_SLICE_X3Y59_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y59_SLICE_X3Y59_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y59_SLICE_X3Y59_CO5),
.O6(CLBLM_R_X3Y59_SLICE_X3Y59_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X3Y59_SLICE_X3Y59_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y59_SLICE_X3Y59_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y59_SLICE_X3Y59_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X3Y59_SLICE_X3Y59_BO5),
.O6(CLBLM_R_X3Y59_SLICE_X3Y59_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X3Y59_SLICE_X3Y59_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y59_SLICE_X3Y59_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y59_SLICE_X3Y59_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X3Y59_SLICE_X3Y59_AO5),
.O6(CLBLM_R_X3Y59_SLICE_X3Y59_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y60_SLICE_X2Y60_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y60_SLICE_X2Y60_DO5),
.O6(CLBLM_R_X3Y60_SLICE_X2Y60_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y60_SLICE_X2Y60_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y60_SLICE_X2Y60_CO5),
.O6(CLBLM_R_X3Y60_SLICE_X2Y60_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y60_SLICE_X2Y60_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y60_SLICE_X2Y60_BO5),
.O6(CLBLM_R_X3Y60_SLICE_X2Y60_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y60_SLICE_X2Y60_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y60_SLICE_X2Y60_AO5),
.O6(CLBLM_R_X3Y60_SLICE_X2Y60_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y60_SLICE_X3Y60_B5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y60_SLICE_X3Y60_BO5),
.Q(CLBLM_R_X3Y60_SLICE_X3Y60_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y60_SLICE_X3Y60_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O),
.CE(1'b1),
.D(CLBLM_R_X3Y60_SLICE_X3Y60_B_XOR),
.Q(CLBLM_R_X3Y60_SLICE_X3Y60_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y60_SLICE_X3Y60_CARRY4 (
.CI(CLBLM_R_X3Y59_SLICE_X3Y59_COUT),
.CO({CLBLM_R_X3Y60_SLICE_X3Y60_COUT, CLBLM_R_X3Y60_SLICE_X3Y60_C_CY, CLBLM_R_X3Y60_SLICE_X3Y60_B_CY, CLBLM_R_X3Y60_SLICE_X3Y60_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X3Y60_SLICE_X3Y60_D_XOR, CLBLM_R_X3Y60_SLICE_X3Y60_C_XOR, CLBLM_R_X3Y60_SLICE_X3Y60_B_XOR, CLBLM_R_X3Y60_SLICE_X3Y60_A_XOR}),
.S({CLBLM_R_X3Y60_SLICE_X3Y60_DO6, CLBLM_R_X3Y60_SLICE_X3Y60_CO6, CLBLM_R_X3Y60_SLICE_X3Y60_BO6, CLBLM_R_X3Y60_SLICE_X3Y60_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaa00000000)
  ) CLBLM_R_X3Y60_SLICE_X3Y60_DLUT (
.I0(1'b0),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y60_SLICE_X3Y60_DO5),
.O6(CLBLM_R_X3Y60_SLICE_X3Y60_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLM_R_X3Y60_SLICE_X3Y60_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b0),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y60_SLICE_X3Y60_CO5),
.O6(CLBLM_R_X3Y60_SLICE_X3Y60_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLM_R_X3Y60_SLICE_X3Y60_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y60_SLICE_X3Y60_BQ),
.I2(1'b1),
.I3(CLBLM_R_X3Y60_SLICE_X3Y60_A_XOR),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y60_SLICE_X3Y60_BO5),
.O6(CLBLM_R_X3Y60_SLICE_X3Y60_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X3Y60_SLICE_X3Y60_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y60_SLICE_X3Y60_B5Q),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y60_SLICE_X3Y60_AO5),
.O6(CLBLM_R_X3Y60_SLICE_X3Y60_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y92_SLICE_X66Y92_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y92_SLICE_X66Y92_DO5),
.O6(CLBLM_R_X41Y92_SLICE_X66Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y92_SLICE_X66Y92_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y92_SLICE_X66Y92_CO5),
.O6(CLBLM_R_X41Y92_SLICE_X66Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y92_SLICE_X66Y92_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y92_SLICE_X66Y92_BO5),
.O6(CLBLM_R_X41Y92_SLICE_X66Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y92_SLICE_X66Y92_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y92_SLICE_X66Y92_AO5),
.O6(CLBLM_R_X41Y92_SLICE_X66Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y92_SLICE_X67Y92_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y92_SLICE_X67Y92_BO5),
.Q(CLBLM_R_X41Y92_SLICE_X67Y92_BQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y92_SLICE_X67Y92_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y92_SLICE_X67Y92_C_XOR),
.Q(CLBLM_R_X41Y92_SLICE_X67Y92_CQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y92_SLICE_X67Y92_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y92_SLICE_X67Y92_DO5),
.Q(CLBLM_R_X41Y92_SLICE_X67Y92_DQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X41Y92_SLICE_X67Y92_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X41Y92_SLICE_X67Y92_D_CY, CLBLM_R_X41Y92_SLICE_X67Y92_C_CY, CLBLM_R_X41Y92_SLICE_X67Y92_B_CY, CLBLM_R_X41Y92_SLICE_X67Y92_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({CLBLM_R_X41Y92_SLICE_X67Y92_D_XOR, CLBLM_R_X41Y92_SLICE_X67Y92_C_XOR, CLBLM_R_X41Y92_SLICE_X67Y92_B_XOR, CLBLM_R_X41Y92_SLICE_X67Y92_A_XOR}),
.S({CLBLM_R_X41Y92_SLICE_X67Y92_DO6, CLBLM_R_X41Y92_SLICE_X67Y92_CO6, CLBLM_R_X41Y92_SLICE_X67Y92_BO6, CLBLM_R_X41Y92_SLICE_X67Y92_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacccccccc)
  ) CLBLM_R_X41Y92_SLICE_X67Y92_DLUT (
.I0(CLBLM_R_X41Y94_SLICE_X67Y94_B5Q),
.I1(CLBLM_R_X41Y92_SLICE_X67Y92_B_XOR),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y92_SLICE_X67Y92_DO5),
.O6(CLBLM_R_X41Y92_SLICE_X67Y92_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0000000000)
  ) CLBLM_R_X41Y92_SLICE_X67Y92_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X41Y92_SLICE_X67Y92_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y92_SLICE_X67Y92_CO5),
.O6(CLBLM_R_X41Y92_SLICE_X67Y92_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLM_R_X41Y92_SLICE_X67Y92_BLUT (
.I0(CLBLM_R_X41Y92_SLICE_X67Y92_AO5),
.I1(CLBLM_R_X41Y92_SLICE_X67Y92_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y92_SLICE_X67Y92_BO5),
.O6(CLBLM_R_X41Y92_SLICE_X67Y92_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff000f0f0f0f)
  ) CLBLM_R_X41Y92_SLICE_X67Y92_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X41Y92_SLICE_X67Y92_BQ),
.I3(CLBLM_R_X41Y92_SLICE_X67Y92_AO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y92_SLICE_X67Y92_AO5),
.O6(CLBLM_R_X41Y92_SLICE_X67Y92_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y93_SLICE_X66Y93_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y93_SLICE_X66Y93_DO5),
.O6(CLBLM_R_X41Y93_SLICE_X66Y93_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y93_SLICE_X66Y93_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y93_SLICE_X66Y93_CO5),
.O6(CLBLM_R_X41Y93_SLICE_X66Y93_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y93_SLICE_X66Y93_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y93_SLICE_X66Y93_BO5),
.O6(CLBLM_R_X41Y93_SLICE_X66Y93_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y93_SLICE_X66Y93_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y93_SLICE_X66Y93_AO5),
.O6(CLBLM_R_X41Y93_SLICE_X66Y93_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y93_SLICE_X67Y93_A5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y93_SLICE_X67Y93_AO5),
.Q(CLBLM_R_X41Y93_SLICE_X67Y93_A5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y93_SLICE_X67Y93_B5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y93_SLICE_X67Y93_BO5),
.Q(CLBLM_R_X41Y93_SLICE_X67Y93_B5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y93_SLICE_X67Y93_C5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y93_SLICE_X67Y93_CO5),
.Q(CLBLM_R_X41Y93_SLICE_X67Y93_C5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y93_SLICE_X67Y93_D5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y93_SLICE_X67Y93_DO5),
.Q(CLBLM_R_X41Y93_SLICE_X67Y93_D5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y93_SLICE_X67Y93_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y93_SLICE_X67Y93_A_XOR),
.Q(CLBLM_R_X41Y93_SLICE_X67Y93_AQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y93_SLICE_X67Y93_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y93_SLICE_X67Y93_B_XOR),
.Q(CLBLM_R_X41Y93_SLICE_X67Y93_BQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y93_SLICE_X67Y93_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y93_SLICE_X67Y93_C_XOR),
.Q(CLBLM_R_X41Y93_SLICE_X67Y93_CQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y93_SLICE_X67Y93_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y93_SLICE_X67Y93_D_XOR),
.Q(CLBLM_R_X41Y93_SLICE_X67Y93_DQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X41Y93_SLICE_X67Y93_CARRY4 (
.CI(CLBLM_R_X41Y92_SLICE_X67Y92_COUT),
.CO({CLBLM_R_X41Y93_SLICE_X67Y93_COUT, CLBLM_R_X41Y93_SLICE_X67Y93_C_CY, CLBLM_R_X41Y93_SLICE_X67Y93_B_CY, CLBLM_R_X41Y93_SLICE_X67Y93_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X41Y93_SLICE_X67Y93_D_XOR, CLBLM_R_X41Y93_SLICE_X67Y93_C_XOR, CLBLM_R_X41Y93_SLICE_X67Y93_B_XOR, CLBLM_R_X41Y93_SLICE_X67Y93_A_XOR}),
.S({CLBLM_R_X41Y93_SLICE_X67Y93_DO6, CLBLM_R_X41Y93_SLICE_X67Y93_CO6, CLBLM_R_X41Y93_SLICE_X67Y93_BO6, CLBLM_R_X41Y93_SLICE_X67Y93_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X41Y93_SLICE_X67Y93_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X41Y95_SLICE_X67Y95_B_XOR),
.I2(CLBLM_R_X41Y93_SLICE_X67Y93_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y93_SLICE_X67Y93_DO5),
.O6(CLBLM_R_X41Y93_SLICE_X67Y93_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccff00ff00)
  ) CLBLM_R_X41Y93_SLICE_X67Y93_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X41Y93_SLICE_X67Y93_CQ),
.I2(1'b1),
.I3(CLBLM_R_X41Y95_SLICE_X67Y95_D_XOR),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y93_SLICE_X67Y93_CO5),
.O6(CLBLM_R_X41Y93_SLICE_X67Y93_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLM_R_X41Y93_SLICE_X67Y93_BLUT (
.I0(CLBLM_R_X41Y95_SLICE_X67Y95_C_XOR),
.I1(CLBLM_R_X41Y93_SLICE_X67Y93_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y93_SLICE_X67Y93_BO5),
.O6(CLBLM_R_X41Y93_SLICE_X67Y93_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X41Y93_SLICE_X67Y93_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X41Y93_SLICE_X67Y93_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X41Y95_SLICE_X67Y95_A_XOR),
.I5(1'b1),
.O5(CLBLM_R_X41Y93_SLICE_X67Y93_AO5),
.O6(CLBLM_R_X41Y93_SLICE_X67Y93_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y94_SLICE_X66Y94_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y94_SLICE_X66Y94_DO5),
.O6(CLBLM_R_X41Y94_SLICE_X66Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y94_SLICE_X66Y94_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y94_SLICE_X66Y94_CO5),
.O6(CLBLM_R_X41Y94_SLICE_X66Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y94_SLICE_X66Y94_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y94_SLICE_X66Y94_BO5),
.O6(CLBLM_R_X41Y94_SLICE_X66Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y94_SLICE_X66Y94_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y94_SLICE_X66Y94_AO5),
.O6(CLBLM_R_X41Y94_SLICE_X66Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y94_SLICE_X67Y94_B5_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y94_SLICE_X67Y94_BO5),
.Q(CLBLM_R_X41Y94_SLICE_X67Y94_B5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y94_SLICE_X67Y94_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y94_SLICE_X67Y94_AO5),
.Q(CLBLM_R_X41Y94_SLICE_X67Y94_AQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y94_SLICE_X67Y94_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y94_SLICE_X67Y94_B_XOR),
.Q(CLBLM_R_X41Y94_SLICE_X67Y94_BQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y94_SLICE_X67Y94_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y94_SLICE_X67Y94_CO5),
.Q(CLBLM_R_X41Y94_SLICE_X67Y94_CQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y94_SLICE_X67Y94_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.D(CLBLM_R_X41Y94_SLICE_X67Y94_DO5),
.Q(CLBLM_R_X41Y94_SLICE_X67Y94_DQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X41Y94_SLICE_X67Y94_CARRY4 (
.CI(CLBLM_R_X41Y93_SLICE_X67Y93_COUT),
.CO({CLBLM_R_X41Y94_SLICE_X67Y94_COUT, CLBLM_R_X41Y94_SLICE_X67Y94_C_CY, CLBLM_R_X41Y94_SLICE_X67Y94_B_CY, CLBLM_R_X41Y94_SLICE_X67Y94_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X41Y94_SLICE_X67Y94_D_XOR, CLBLM_R_X41Y94_SLICE_X67Y94_C_XOR, CLBLM_R_X41Y94_SLICE_X67Y94_B_XOR, CLBLM_R_X41Y94_SLICE_X67Y94_A_XOR}),
.S({CLBLM_R_X41Y94_SLICE_X67Y94_DO6, CLBLM_R_X41Y94_SLICE_X67Y94_CO6, CLBLM_R_X41Y94_SLICE_X67Y94_BO6, CLBLM_R_X41Y94_SLICE_X67Y94_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaaaaaaa)
  ) CLBLM_R_X41Y94_SLICE_X67Y94_DLUT (
.I0(CLBLM_R_X41Y94_SLICE_X67Y94_C_XOR),
.I1(1'b1),
.I2(CLBLM_R_X41Y94_SLICE_X67Y94_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y94_SLICE_X67Y94_DO5),
.O6(CLBLM_R_X41Y94_SLICE_X67Y94_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X41Y94_SLICE_X67Y94_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X41Y94_SLICE_X67Y94_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X41Y94_SLICE_X67Y94_A_XOR),
.I5(1'b1),
.O5(CLBLM_R_X41Y94_SLICE_X67Y94_CO5),
.O6(CLBLM_R_X41Y94_SLICE_X67Y94_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLM_R_X41Y94_SLICE_X67Y94_BLUT (
.I0(CLBLM_R_X41Y92_SLICE_X67Y92_D_XOR),
.I1(CLBLM_R_X41Y94_SLICE_X67Y94_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y94_SLICE_X67Y94_BO5),
.O6(CLBLM_R_X41Y94_SLICE_X67Y94_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0f0f0f0)
  ) CLBLM_R_X41Y94_SLICE_X67Y94_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X41Y94_SLICE_X67Y94_CQ),
.I2(CLBLM_R_X41Y94_SLICE_X67Y94_D_XOR),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y94_SLICE_X67Y94_AO5),
.O6(CLBLM_R_X41Y94_SLICE_X67Y94_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y95_SLICE_X66Y95_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y95_SLICE_X66Y95_DO5),
.O6(CLBLM_R_X41Y95_SLICE_X66Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y95_SLICE_X66Y95_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y95_SLICE_X66Y95_CO5),
.O6(CLBLM_R_X41Y95_SLICE_X66Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y95_SLICE_X66Y95_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y95_SLICE_X66Y95_BO5),
.O6(CLBLM_R_X41Y95_SLICE_X66Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y95_SLICE_X66Y95_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y95_SLICE_X66Y95_AO5),
.O6(CLBLM_R_X41Y95_SLICE_X66Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y95_SLICE_X67Y95_A_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y95_SLICE_X67Y95_AO5),
.Q(CLBLM_R_X41Y95_SLICE_X67Y95_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y95_SLICE_X67Y95_B_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y95_SLICE_X67Y95_BO5),
.Q(CLBLM_R_X41Y95_SLICE_X67Y95_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y95_SLICE_X67Y95_C_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y95_SLICE_X67Y95_CO5),
.Q(CLBLM_R_X41Y95_SLICE_X67Y95_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y95_SLICE_X67Y95_D_FDRE (
.C(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y95_SLICE_X67Y95_DO5),
.Q(CLBLM_R_X41Y95_SLICE_X67Y95_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X41Y95_SLICE_X67Y95_CARRY4 (
.CI(CLBLM_R_X41Y94_SLICE_X67Y94_COUT),
.CO({CLBLM_R_X41Y95_SLICE_X67Y95_COUT, CLBLM_R_X41Y95_SLICE_X67Y95_C_CY, CLBLM_R_X41Y95_SLICE_X67Y95_B_CY, CLBLM_R_X41Y95_SLICE_X67Y95_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X41Y95_SLICE_X67Y95_D_XOR, CLBLM_R_X41Y95_SLICE_X67Y95_C_XOR, CLBLM_R_X41Y95_SLICE_X67Y95_B_XOR, CLBLM_R_X41Y95_SLICE_X67Y95_A_XOR}),
.S({CLBLM_R_X41Y95_SLICE_X67Y95_DO6, CLBLM_R_X41Y95_SLICE_X67Y95_CO6, CLBLM_R_X41Y95_SLICE_X67Y95_BO6, CLBLM_R_X41Y95_SLICE_X67Y95_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00ffff0000)
  ) CLBLM_R_X41Y95_SLICE_X67Y95_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X41Y93_SLICE_X67Y93_C5Q),
.I4(CLBLM_R_X41Y94_SLICE_X67Y94_AQ),
.I5(1'b1),
.O5(CLBLM_R_X41Y95_SLICE_X67Y95_DO5),
.O6(CLBLM_R_X41Y95_SLICE_X67Y95_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacccccccc)
  ) CLBLM_R_X41Y95_SLICE_X67Y95_CLUT (
.I0(CLBLM_R_X41Y93_SLICE_X67Y93_B5Q),
.I1(CLBLM_R_X41Y93_SLICE_X67Y93_A5Q),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y95_SLICE_X67Y95_CO5),
.O6(CLBLM_R_X41Y95_SLICE_X67Y95_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaf0f0f0f0)
  ) CLBLM_R_X41Y95_SLICE_X67Y95_BLUT (
.I0(CLBLM_R_X41Y93_SLICE_X67Y93_D5Q),
.I1(1'b1),
.I2(CLBLM_R_X41Y93_SLICE_X67Y93_B5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y95_SLICE_X67Y95_BO5),
.O6(CLBLM_R_X41Y95_SLICE_X67Y95_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaaaaaaa)
  ) CLBLM_R_X41Y95_SLICE_X67Y95_ALUT (
.I0(CLBLM_R_X41Y93_SLICE_X67Y93_D5Q),
.I1(1'b1),
.I2(CLBLM_R_X41Y93_SLICE_X67Y93_A5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y95_SLICE_X67Y95_AO5),
.O6(CLBLM_R_X41Y95_SLICE_X67Y95_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y100_SLICE_X66Y100_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y100_SLICE_X66Y100_DO5),
.O6(CLBLM_R_X41Y100_SLICE_X66Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y100_SLICE_X66Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y100_SLICE_X66Y100_CO5),
.O6(CLBLM_R_X41Y100_SLICE_X66Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y100_SLICE_X66Y100_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y100_SLICE_X66Y100_BO5),
.O6(CLBLM_R_X41Y100_SLICE_X66Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y100_SLICE_X66Y100_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y100_SLICE_X66Y100_AO5),
.O6(CLBLM_R_X41Y100_SLICE_X66Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y100_SLICE_X67Y100_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y100_SLICE_X67Y100_AO5),
.Q(CLBLM_R_X41Y100_SLICE_X67Y100_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y100_SLICE_X67Y100_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y100_SLICE_X67Y100_CO5),
.Q(CLBLM_R_X41Y100_SLICE_X67Y100_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y100_SLICE_X67Y100_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y100_SLICE_X67Y100_DO5),
.Q(CLBLM_R_X41Y100_SLICE_X67Y100_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y100_SLICE_X67Y100_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y92_SLICE_X67Y92_BQ),
.Q(CLBLM_R_X41Y100_SLICE_X67Y100_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y100_SLICE_X67Y100_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y94_SLICE_X67Y94_B5Q),
.Q(CLBLM_R_X41Y100_SLICE_X67Y100_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y100_SLICE_X67Y100_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y93_SLICE_X67Y93_CQ),
.Q(CLBLM_R_X41Y100_SLICE_X67Y100_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y100_SLICE_X67Y100_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y92_SLICE_X67Y92_CQ),
.Q(CLBLM_R_X41Y100_SLICE_X67Y100_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaaaaaa)
  ) CLBLM_R_X41Y100_SLICE_X67Y100_DLUT (
.I0(CLBLM_R_X41Y92_SLICE_X67Y92_DQ),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y100_SLICE_X67Y100_DO5),
.O6(CLBLM_R_X41Y100_SLICE_X67Y100_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f0f0f0f0)
  ) CLBLM_R_X41Y100_SLICE_X67Y100_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X41Y93_SLICE_X67Y93_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y100_SLICE_X67Y100_CO5),
.O6(CLBLM_R_X41Y100_SLICE_X67Y100_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000e400e400)
  ) CLBLM_R_X41Y100_SLICE_X67Y100_BLUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I1(CLBLM_R_X41Y107_SLICE_X66Y107_DO6),
.I2(CLBLM_R_X41Y103_SLICE_X67Y103_BO6),
.I3(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y100_SLICE_X67Y100_BO5),
.O6(CLBLM_R_X41Y100_SLICE_X67Y100_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLM_R_X41Y100_SLICE_X67Y100_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X41Y93_SLICE_X67Y93_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y100_SLICE_X67Y100_AO5),
.O6(CLBLM_R_X41Y100_SLICE_X67Y100_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000ff0000)
  ) CLBLM_R_X41Y101_SLICE_X66Y101_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X41Y110_SLICE_X66Y110_DO5),
.I4(CLBLL_L_X42Y110_SLICE_X68Y110_BO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y101_SLICE_X66Y101_DO5),
.O6(CLBLM_R_X41Y101_SLICE_X66Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000045004000)
  ) CLBLM_R_X41Y101_SLICE_X66Y101_CLUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I1(CLBLM_R_X41Y105_SLICE_X66Y105_CO6),
.I2(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I3(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I4(CLBLM_R_X41Y105_SLICE_X67Y105_AO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y101_SLICE_X66Y101_CO5),
.O6(CLBLM_R_X41Y101_SLICE_X66Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000005d7f)
  ) CLBLM_R_X41Y101_SLICE_X66Y101_BLUT (
.I0(CLBLM_R_X41Y105_SLICE_X67Y105_CO6),
.I1(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I2(CLBLL_L_X42Y107_SLICE_X68Y107_AO6),
.I3(CLBLM_R_X41Y104_SLICE_X66Y104_DO6),
.I4(CLBLM_R_X41Y101_SLICE_X66Y101_CO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y101_SLICE_X66Y101_BO5),
.O6(CLBLM_R_X41Y101_SLICE_X66Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y101_SLICE_X66Y101_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y101_SLICE_X66Y101_AO5),
.O6(CLBLM_R_X41Y101_SLICE_X66Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y101_SLICE_X67Y101_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y102_SLICE_X67Y102_DO5),
.D(CLBLM_R_X41Y101_SLICE_X67Y101_AO6),
.Q(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y101_SLICE_X67Y101_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y102_SLICE_X67Y102_DO5),
.D(CLBLM_R_X41Y101_SLICE_X67Y101_DO5),
.Q(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y101_SLICE_X67Y101_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y102_SLICE_X67Y102_DO5),
.D(CLBLM_R_X41Y101_SLICE_X67Y101_CO6),
.Q(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h88008800ffff0000)
  ) CLBLM_R_X41Y101_SLICE_X67Y101_DLUT (
.I0(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I1(CLBLL_L_X42Y105_SLICE_X69Y105_DO5),
.I2(1'b1),
.I3(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I4(CLBLM_R_X41Y101_SLICE_X67Y101_AO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y101_SLICE_X67Y101_DO5),
.O6(CLBLM_R_X41Y101_SLICE_X67Y101_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0c0c0c000000000)
  ) CLBLM_R_X41Y101_SLICE_X67Y101_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y110_SLICE_X68Y110_BO5),
.I2(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y101_SLICE_X67Y101_CO5),
.O6(CLBLM_R_X41Y101_SLICE_X67Y101_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000020222000)
  ) CLBLM_R_X41Y101_SLICE_X67Y101_BLUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I1(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I2(CLBLL_L_X42Y107_SLICE_X68Y107_AO6),
.I3(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I4(CLBLM_R_X41Y104_SLICE_X66Y104_DO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y101_SLICE_X67Y101_BO5),
.O6(CLBLM_R_X41Y101_SLICE_X67Y101_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00f000f000)
  ) CLBLM_R_X41Y101_SLICE_X67Y101_ALUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I1(1'b1),
.I2(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I3(CLBLL_L_X42Y110_SLICE_X68Y110_BO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y101_SLICE_X67Y101_AO5),
.O6(CLBLM_R_X41Y101_SLICE_X67Y101_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y102_SLICE_X66Y102_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLM_R_X41Y102_SLICE_X66Y102_DO5),
.Q(CLBLM_R_X41Y102_SLICE_X66Y102_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000077007000)
  ) CLBLM_R_X41Y102_SLICE_X66Y102_DLUT (
.I0(CLBLL_L_X42Y103_SLICE_X68Y103_CO6),
.I1(CLBLM_R_X41Y108_SLICE_X67Y108_BO6),
.I2(CLBLL_L_X42Y97_SLICE_X69Y97_C5Q),
.I3(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I4(CLBLM_R_X41Y102_SLICE_X66Y102_BQ),
.I5(1'b1),
.O5(CLBLM_R_X41Y102_SLICE_X66Y102_DO5),
.O6(CLBLM_R_X41Y102_SLICE_X66Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000033330f0a0f0a)
  ) CLBLM_R_X41Y102_SLICE_X66Y102_CLUT (
.I0(CLBLL_L_X42Y103_SLICE_X68Y103_CO6),
.I1(CLBLM_R_X41Y108_SLICE_X67Y108_BO6),
.I2(CLBLM_R_X41Y115_SLICE_X66Y115_DO6),
.I3(CLBLM_R_X41Y102_SLICE_X66Y102_CO6),
.I4(CLBLM_R_X41Y107_SLICE_X66Y107_AO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y102_SLICE_X66Y102_CO5),
.O6(CLBLM_R_X41Y102_SLICE_X66Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ccc0ccc0)
  ) CLBLM_R_X41Y102_SLICE_X66Y102_BLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y102_SLICE_X68Y102_AO6),
.I2(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.I3(CLBLM_R_X41Y105_SLICE_X67Y105_CO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y102_SLICE_X66Y102_BO5),
.O6(CLBLM_R_X41Y102_SLICE_X66Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f00002020aaa)
  ) CLBLM_R_X41Y102_SLICE_X66Y102_ALUT (
.I0(CLBLM_R_X41Y102_SLICE_X66Y102_CO5),
.I1(CLBLL_L_X42Y109_SLICE_X69Y109_CO6),
.I2(CLBLM_R_X41Y109_SLICE_X67Y109_CO6),
.I3(CLBLM_R_X41Y102_SLICE_X66Y102_BO5),
.I4(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I5(1'b1),
.O5(CLBLM_R_X41Y102_SLICE_X66Y102_AO5),
.O6(CLBLM_R_X41Y102_SLICE_X66Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y102_SLICE_X67Y102_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y102_SLICE_X67Y102_AO5),
.D(CLBLM_R_X41Y102_SLICE_X67Y102_CO5),
.Q(CLBLM_R_X41Y102_SLICE_X67Y102_C5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000010)
  ) CLBLM_R_X41Y102_SLICE_X67Y102_DLUT (
.I0(CLBLM_R_X41Y109_SLICE_X66Y109_BO5),
.I1(CLBLM_R_X41Y108_SLICE_X67Y108_BO6),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(CLBLL_L_X42Y109_SLICE_X69Y109_BO5),
.I4(CLBLM_R_X41Y102_SLICE_X67Y102_BO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y102_SLICE_X67Y102_DO5),
.O6(CLBLM_R_X41Y102_SLICE_X67Y102_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000a4e0a4e)
  ) CLBLM_R_X41Y102_SLICE_X67Y102_CLUT (
.I0(CLBLL_L_X42Y109_SLICE_X69Y109_CO6),
.I1(CLBLM_R_X41Y109_SLICE_X67Y109_CO6),
.I2(CLBLL_L_X42Y103_SLICE_X68Y103_CO6),
.I3(CLBLM_R_X41Y102_SLICE_X66Y102_BO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y102_SLICE_X67Y102_CO5),
.O6(CLBLM_R_X41Y102_SLICE_X67Y102_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000c0ff)
  ) CLBLM_R_X41Y102_SLICE_X67Y102_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X41Y102_SLICE_X66Y102_BO5),
.I2(CLBLL_L_X42Y102_SLICE_X68Y102_CO6),
.I3(CLBLL_L_X42Y102_SLICE_X68Y102_DO6),
.I4(CLBLL_L_X42Y103_SLICE_X68Y103_CO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y102_SLICE_X67Y102_BO5),
.O6(CLBLM_R_X41Y102_SLICE_X67Y102_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000550055)
  ) CLBLM_R_X41Y102_SLICE_X67Y102_ALUT (
.I0(CLBLM_R_X41Y115_SLICE_X66Y115_DO6),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X41Y109_SLICE_X66Y109_BO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y102_SLICE_X67Y102_AO5),
.O6(CLBLM_R_X41Y102_SLICE_X67Y102_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y103_SLICE_X66Y103_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y103_SLICE_X66Y103_DO5),
.O6(CLBLM_R_X41Y103_SLICE_X66Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000a022f577)
  ) CLBLM_R_X41Y103_SLICE_X66Y103_CLUT (
.I0(CLBLL_L_X42Y109_SLICE_X69Y109_BO5),
.I1(CLBLM_R_X41Y109_SLICE_X67Y109_BO5),
.I2(CLBLM_R_X41Y104_SLICE_X67Y104_C5Q),
.I3(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I4(CLBLM_R_X41Y103_SLICE_X66Y103_BO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y103_SLICE_X66Y103_CO5),
.O6(CLBLM_R_X41Y103_SLICE_X66Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000007770777)
  ) CLBLM_R_X41Y103_SLICE_X66Y103_BLUT (
.I0(CLBLL_L_X42Y110_SLICE_X68Y110_AO5),
.I1(CLBLM_R_X41Y114_SLICE_X67Y114_A5Q),
.I2(CLBLM_R_X41Y111_SLICE_X66Y111_DQ),
.I3(CLBLM_R_X41Y109_SLICE_X67Y109_CO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y103_SLICE_X66Y103_BO5),
.O6(CLBLM_R_X41Y103_SLICE_X66Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X41Y103_SLICE_X66Y103_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y103_SLICE_X66Y103_AO5),
.O6(CLBLM_R_X41Y103_SLICE_X66Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y103_SLICE_X67Y103_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y110_SLICE_X68Y110_BO6),
.D(CLBLM_R_X41Y103_SLICE_X67Y103_DO5),
.Q(CLBLM_R_X41Y103_SLICE_X67Y103_D5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff80ff)
  ) CLBLM_R_X41Y103_SLICE_X67Y103_DLUT (
.I0(CLBLL_L_X42Y109_SLICE_X69Y109_BO5),
.I1(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I2(CLBLM_R_X41Y103_SLICE_X67Y103_D5Q),
.I3(CLBLM_R_X41Y116_SLICE_X67Y116_DO5),
.I4(CLBLM_R_X41Y103_SLICE_X67Y103_AO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y103_SLICE_X67Y103_DO5),
.O6(CLBLM_R_X41Y103_SLICE_X67Y103_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000aaaafc30)
  ) CLBLM_R_X41Y103_SLICE_X67Y103_CLUT (
.I0(CLBLM_R_X41Y106_SLICE_X66Y106_BO6),
.I1(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I2(CLBLM_R_X41Y105_SLICE_X67Y105_AO6),
.I3(CLBLM_R_X41Y105_SLICE_X66Y105_CO6),
.I4(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I5(1'b1),
.O5(CLBLM_R_X41Y103_SLICE_X67Y103_CO5),
.O6(CLBLM_R_X41Y103_SLICE_X67Y103_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hd0dff0ff808ff0ff)
  ) CLBLM_R_X41Y103_SLICE_X67Y103_BLUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I1(CLBLL_L_X42Y106_SLICE_X68Y106_CO5),
.I2(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I3(CLBLL_L_X42Y105_SLICE_X69Y105_BO5),
.I4(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I5(CLBLL_L_X42Y101_SLICE_X69Y101_DO6),
.O5(CLBLM_R_X41Y103_SLICE_X67Y103_BO5),
.O6(CLBLM_R_X41Y103_SLICE_X67Y103_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h020a222a00082028)
  ) CLBLM_R_X41Y103_SLICE_X67Y103_ALUT (
.I0(CLBLM_R_X41Y107_SLICE_X67Y107_BO6),
.I1(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I2(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.I3(CLBLM_R_X41Y107_SLICE_X66Y107_DO6),
.I4(CLBLM_R_X41Y103_SLICE_X67Y103_BO6),
.I5(CLBLM_R_X41Y103_SLICE_X67Y103_CO5),
.O5(CLBLM_R_X41Y103_SLICE_X67Y103_AO5),
.O6(CLBLM_R_X41Y103_SLICE_X67Y103_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y104_SLICE_X66Y104_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y101_SLICE_X66Y101_DO5),
.D(CLBLM_R_X41Y104_SLICE_X66Y104_AO6),
.Q(CLBLM_R_X41Y104_SLICE_X66Y104_D5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hc044c04400000000)
  ) CLBLM_R_X41Y104_SLICE_X66Y104_DLUT (
.I0(CLBLL_L_X42Y102_SLICE_X69Y102_BO5),
.I1(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I2(CLBLM_R_X41Y100_SLICE_X67Y100_DQ),
.I3(CLBLL_L_X42Y107_SLICE_X68Y107_BO5),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y104_SLICE_X66Y104_DO5),
.O6(CLBLM_R_X41Y104_SLICE_X66Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h777700000f000f00)
  ) CLBLM_R_X41Y104_SLICE_X66Y104_CLUT (
.I0(CLBLM_R_X41Y109_SLICE_X67Y109_DO6),
.I1(CLBLL_L_X42Y109_SLICE_X69Y109_BO5),
.I2(CLBLM_R_X41Y105_SLICE_X66Y105_AO6),
.I3(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I4(CLBLM_R_X41Y109_SLICE_X67Y109_AO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y104_SLICE_X66Y104_CO5),
.O6(CLBLM_R_X41Y104_SLICE_X66Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000001333133)
  ) CLBLM_R_X41Y104_SLICE_X66Y104_BLUT (
.I0(CLBLL_L_X42Y107_SLICE_X68Y107_CO6),
.I1(CLBLM_R_X41Y105_SLICE_X67Y105_CO5),
.I2(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I3(CLBLM_R_X41Y105_SLICE_X67Y105_CO6),
.I4(CLBLM_R_X41Y104_SLICE_X66Y104_DO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y104_SLICE_X66Y104_BO5),
.O6(CLBLM_R_X41Y104_SLICE_X66Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hbb3bbb3bbb33bb3b)
  ) CLBLM_R_X41Y104_SLICE_X66Y104_ALUT (
.I0(CLBLM_R_X41Y107_SLICE_X67Y107_BO6),
.I1(CLBLM_R_X41Y104_SLICE_X66Y104_CO6),
.I2(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.I3(CLBLL_L_X42Y104_SLICE_X68Y104_CO6),
.I4(CLBLM_R_X41Y104_SLICE_X66Y104_BO5),
.I5(CLBLM_R_X41Y104_SLICE_X66Y104_CO5),
.O5(CLBLM_R_X41Y104_SLICE_X66Y104_AO5),
.O6(CLBLM_R_X41Y104_SLICE_X66Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y104_SLICE_X67Y104_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y110_SLICE_X68Y110_BO6),
.D(CLBLM_R_X41Y104_SLICE_X67Y104_AO6),
.Q(CLBLM_R_X41Y104_SLICE_X67Y104_C5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h3300330044444444)
  ) CLBLM_R_X41Y104_SLICE_X67Y104_DLUT (
.I0(CLBLL_L_X42Y105_SLICE_X68Y105_CO5),
.I1(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I2(1'b1),
.I3(CLBLL_L_X42Y105_SLICE_X68Y105_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y104_SLICE_X67Y104_DO5),
.O6(CLBLM_R_X41Y104_SLICE_X67Y104_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hc0ccc00000000000)
  ) CLBLM_R_X41Y104_SLICE_X67Y104_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X41Y105_SLICE_X67Y105_CO6),
.I2(CLBLM_R_X41Y105_SLICE_X67Y105_AO6),
.I3(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I4(CLBLL_L_X42Y107_SLICE_X68Y107_AO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y104_SLICE_X67Y104_CO5),
.O6(CLBLM_R_X41Y104_SLICE_X67Y104_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000f0f0e0c)
  ) CLBLM_R_X41Y104_SLICE_X67Y104_BLUT (
.I0(CLBLL_L_X42Y105_SLICE_X68Y105_CO6),
.I1(CLBLL_L_X42Y103_SLICE_X68Y103_AO6),
.I2(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.I3(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I4(CLBLM_R_X41Y104_SLICE_X67Y104_CO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y104_SLICE_X67Y104_BO5),
.O6(CLBLM_R_X41Y104_SLICE_X67Y104_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffffaaaaffff0020)
  ) CLBLM_R_X41Y104_SLICE_X67Y104_ALUT (
.I0(CLBLM_R_X41Y107_SLICE_X67Y107_BO6),
.I1(CLBLM_R_X41Y104_SLICE_X67Y104_DO5),
.I2(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.I3(CLBLM_R_X41Y104_SLICE_X67Y104_DO6),
.I4(CLBLM_R_X41Y103_SLICE_X66Y103_CO5),
.I5(CLBLM_R_X41Y104_SLICE_X67Y104_BO5),
.O5(CLBLM_R_X41Y104_SLICE_X67Y104_AO5),
.O6(CLBLM_R_X41Y104_SLICE_X67Y104_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y105_SLICE_X66Y105_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y110_SLICE_X68Y110_BO6),
.D(CLBLM_R_X41Y105_SLICE_X66Y105_DO6),
.Q(CLBLM_R_X41Y105_SLICE_X66Y105_DQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h33333333f3f3f373)
  ) CLBLM_R_X41Y105_SLICE_X66Y105_DLUT (
.I0(CLBLL_L_X42Y106_SLICE_X69Y106_BO5),
.I1(CLBLM_R_X41Y111_SLICE_X67Y111_DO5),
.I2(CLBLM_R_X41Y107_SLICE_X67Y107_BO6),
.I3(CLBLM_R_X41Y101_SLICE_X67Y101_BO5),
.I4(CLBLM_R_X41Y105_SLICE_X66Y105_BO6),
.I5(CLBLM_R_X41Y100_SLICE_X67Y100_BO5),
.O5(CLBLM_R_X41Y105_SLICE_X66Y105_DO5),
.O6(CLBLM_R_X41Y105_SLICE_X66Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h88888888aaa00a00)
  ) CLBLM_R_X41Y105_SLICE_X66Y105_CLUT (
.I0(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I1(CLBLM_R_X41Y100_SLICE_X67Y100_C5Q),
.I2(CLBLM_R_X41Y108_SLICE_X66Y108_CO6),
.I3(CLBLL_L_X42Y108_SLICE_X69Y108_BO5),
.I4(CLBLL_L_X42Y102_SLICE_X69Y102_C5Q),
.I5(CLBLL_L_X42Y107_SLICE_X68Y107_BO5),
.O5(CLBLM_R_X41Y105_SLICE_X66Y105_CO5),
.O6(CLBLM_R_X41Y105_SLICE_X66Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0a0e0e050004040)
  ) CLBLM_R_X41Y105_SLICE_X66Y105_BLUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I1(CLBLM_R_X41Y105_SLICE_X67Y105_AO6),
.I2(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I3(CLBLM_R_X41Y105_SLICE_X66Y105_CO6),
.I4(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I5(CLBLM_R_X41Y106_SLICE_X66Y106_BO6),
.O5(CLBLM_R_X41Y105_SLICE_X66Y105_BO5),
.O6(CLBLM_R_X41Y105_SLICE_X66Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0c040f07fcf4fff7)
  ) CLBLM_R_X41Y105_SLICE_X66Y105_ALUT (
.I0(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I1(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I2(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I3(CLBLM_R_X41Y106_SLICE_X66Y106_CO6),
.I4(CLBLM_R_X41Y105_SLICE_X66Y105_CO6),
.I5(CLBLM_R_X41Y106_SLICE_X66Y106_AO6),
.O5(CLBLM_R_X41Y105_SLICE_X66Y105_AO5),
.O6(CLBLM_R_X41Y105_SLICE_X66Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000a2aaaaaa)
  ) CLBLM_R_X41Y105_SLICE_X67Y105_DLUT (
.I0(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I1(CLBLM_R_X41Y109_SLICE_X66Y109_BO6),
.I2(CLBLM_R_X41Y100_SLICE_X67Y100_A5Q),
.I3(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I4(CLBLL_L_X42Y109_SLICE_X69Y109_DQ),
.I5(1'b1),
.O5(CLBLM_R_X41Y105_SLICE_X67Y105_DO5),
.O6(CLBLM_R_X41Y105_SLICE_X67Y105_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003332001000)
  ) CLBLM_R_X41Y105_SLICE_X67Y105_CLUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I1(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I2(CLBLL_L_X42Y107_SLICE_X68Y107_AO6),
.I3(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I4(CLBLM_R_X41Y105_SLICE_X67Y105_AO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y105_SLICE_X67Y105_CO5),
.O6(CLBLM_R_X41Y105_SLICE_X67Y105_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000331333b3)
  ) CLBLM_R_X41Y105_SLICE_X67Y105_BLUT (
.I0(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I1(CLBLL_L_X42Y107_SLICE_X69Y107_CQ),
.I2(CLBLM_R_X41Y108_SLICE_X67Y108_BO6),
.I3(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I4(CLBLL_L_X42Y108_SLICE_X69Y108_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X41Y105_SLICE_X67Y105_BO5),
.O6(CLBLM_R_X41Y105_SLICE_X67Y105_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hc8c08800c8c0cccc)
  ) CLBLM_R_X41Y105_SLICE_X67Y105_ALUT (
.I0(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I1(CLBLM_R_X41Y105_SLICE_X67Y105_DO5),
.I2(CLBLL_L_X42Y107_SLICE_X69Y107_DQ),
.I3(CLBLM_R_X41Y107_SLICE_X66Y107_AO6),
.I4(CLBLM_R_X41Y108_SLICE_X66Y108_CO6),
.I5(CLBLM_R_X41Y105_SLICE_X67Y105_BO5),
.O5(CLBLM_R_X41Y105_SLICE_X67Y105_AO5),
.O6(CLBLM_R_X41Y105_SLICE_X67Y105_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000050c55cc)
  ) CLBLM_R_X41Y106_SLICE_X66Y106_DLUT (
.I0(CLBLL_L_X42Y107_SLICE_X69Y107_BQ),
.I1(CLBLL_L_X42Y108_SLICE_X68Y108_BO5),
.I2(CLBLM_R_X41Y107_SLICE_X66Y107_AO6),
.I3(CLBLM_R_X41Y108_SLICE_X66Y108_CO6),
.I4(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y106_SLICE_X66Y106_DO5),
.O6(CLBLM_R_X41Y106_SLICE_X66Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h27770fff227200f0)
  ) CLBLM_R_X41Y106_SLICE_X66Y106_CLUT (
.I0(CLBLM_R_X41Y107_SLICE_X66Y107_AO6),
.I1(CLBLM_R_X41Y100_SLICE_X67Y100_CQ),
.I2(CLBLM_R_X41Y108_SLICE_X66Y108_CO6),
.I3(CLBLL_L_X42Y107_SLICE_X69Y107_D5Q),
.I4(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I5(CLBLL_L_X42Y106_SLICE_X68Y106_BO5),
.O5(CLBLM_R_X41Y106_SLICE_X66Y106_CO5),
.O6(CLBLM_R_X41Y106_SLICE_X66Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h2000202070507070)
  ) CLBLM_R_X41Y106_SLICE_X66Y106_BLUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I1(CLBLM_R_X41Y106_SLICE_X66Y106_DO5),
.I2(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I3(CLBLM_R_X41Y106_SLICE_X67Y106_BQ),
.I4(CLBLL_L_X42Y107_SLICE_X68Y107_BO5),
.I5(CLBLM_R_X41Y106_SLICE_X66Y106_CO6),
.O5(CLBLM_R_X41Y106_SLICE_X66Y106_BO5),
.O6(CLBLM_R_X41Y106_SLICE_X66Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000b00f000fb00)
  ) CLBLM_R_X41Y106_SLICE_X66Y106_ALUT (
.I0(CLBLM_R_X41Y106_SLICE_X67Y106_BQ),
.I1(CLBLL_L_X42Y107_SLICE_X68Y107_BO5),
.I2(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I3(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I4(CLBLM_R_X41Y106_SLICE_X66Y106_DO5),
.I5(CLBLM_R_X41Y107_SLICE_X66Y107_CO6),
.O5(CLBLM_R_X41Y106_SLICE_X66Y106_AO5),
.O6(CLBLM_R_X41Y106_SLICE_X66Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y106_SLICE_X67Y106_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y106_SLICE_X67Y106_AO5),
.Q(CLBLM_R_X41Y106_SLICE_X67Y106_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y106_SLICE_X67Y106_C5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y106_SLICE_X67Y106_CO5),
.Q(CLBLM_R_X41Y106_SLICE_X67Y106_C5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y106_SLICE_X67Y106_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y114_SLICE_X66Y114_D5Q),
.Q(CLBLM_R_X41Y106_SLICE_X67Y106_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y106_SLICE_X67Y106_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y93_SLICE_X67Y93_DQ),
.Q(CLBLM_R_X41Y106_SLICE_X67Y106_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y106_SLICE_X67Y106_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y94_SLICE_X67Y94_DQ),
.Q(CLBLM_R_X41Y106_SLICE_X67Y106_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000a0a08800)
  ) CLBLM_R_X41Y106_SLICE_X67Y106_DLUT (
.I0(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I1(CLBLM_R_X41Y108_SLICE_X67Y108_CO6),
.I2(CLBLM_R_X41Y106_SLICE_X67Y106_CQ),
.I3(CLBLL_L_X42Y111_SLICE_X69Y111_DQ),
.I4(CLBLL_L_X42Y106_SLICE_X69Y106_CO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y106_SLICE_X67Y106_DO5),
.O6(CLBLM_R_X41Y106_SLICE_X67Y106_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff00ff00)
  ) CLBLM_R_X41Y106_SLICE_X67Y106_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X41Y94_SLICE_X67Y94_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y106_SLICE_X67Y106_CO5),
.O6(CLBLM_R_X41Y106_SLICE_X67Y106_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'haa0aa000aa00aa00)
  ) CLBLM_R_X41Y106_SLICE_X67Y106_BLUT (
.I0(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I1(1'b1),
.I2(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I3(CLBLM_R_X41Y106_SLICE_X67Y106_DO5),
.I4(CLBLM_R_X41Y107_SLICE_X66Y107_BO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y106_SLICE_X67Y106_BO5),
.O6(CLBLM_R_X41Y106_SLICE_X67Y106_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cccccccc)
  ) CLBLM_R_X41Y106_SLICE_X67Y106_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X41Y94_SLICE_X67Y94_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y106_SLICE_X67Y106_AO5),
.O6(CLBLM_R_X41Y106_SLICE_X67Y106_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0500af220555af77)
  ) CLBLM_R_X41Y107_SLICE_X66Y107_DLUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I1(CLBLM_R_X41Y106_SLICE_X67Y106_BO5),
.I2(CLBLM_R_X41Y107_SLICE_X66Y107_BO6),
.I3(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I4(CLBLM_R_X41Y101_SLICE_X67Y101_DO6),
.I5(CLBLM_R_X41Y107_SLICE_X67Y107_BO5),
.O5(CLBLM_R_X41Y107_SLICE_X66Y107_DO5),
.O6(CLBLM_R_X41Y107_SLICE_X66Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h002ac0ea153fd5ff)
  ) CLBLM_R_X41Y107_SLICE_X66Y107_CLUT (
.I0(CLBLM_R_X41Y108_SLICE_X66Y108_CO6),
.I1(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I2(CLBLM_R_X41Y107_SLICE_X66Y107_AO6),
.I3(CLBLL_L_X42Y107_SLICE_X69Y107_B5Q),
.I4(CLBLM_R_X41Y106_SLICE_X67Y106_A5Q),
.I5(CLBLL_L_X42Y108_SLICE_X68Y108_DO5),
.O5(CLBLM_R_X41Y107_SLICE_X66Y107_CO5),
.O6(CLBLM_R_X41Y107_SLICE_X66Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hfaaafccc00000000)
  ) CLBLM_R_X41Y107_SLICE_X66Y107_BLUT (
.I0(CLBLL_L_X42Y68_SLICE_X68Y68_BQ),
.I1(CLBLL_L_X42Y108_SLICE_X68Y108_AO5),
.I2(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I3(CLBLM_R_X41Y107_SLICE_X66Y107_AO6),
.I4(CLBLM_R_X41Y108_SLICE_X66Y108_CO6),
.I5(CLBLL_L_X42Y107_SLICE_X68Y107_BO6),
.O5(CLBLM_R_X41Y107_SLICE_X66Y107_BO5),
.O6(CLBLM_R_X41Y107_SLICE_X66Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100000000000000)
  ) CLBLM_R_X41Y107_SLICE_X66Y107_ALUT (
.I0(CLBLM_R_X41Y108_SLICE_X66Y108_D5Q),
.I1(CLBLM_R_X41Y109_SLICE_X66Y109_AQ),
.I2(CLBLL_L_X42Y109_SLICE_X68Y109_DQ),
.I3(CLBLM_R_X41Y108_SLICE_X67Y108_CO5),
.I4(CLBLL_L_X42Y106_SLICE_X69Y106_CO6),
.I5(CLBLM_R_X41Y108_SLICE_X67Y108_DO6),
.O5(CLBLM_R_X41Y107_SLICE_X66Y107_AO5),
.O6(CLBLM_R_X41Y107_SLICE_X66Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y107_SLICE_X67Y107_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y110_SLICE_X68Y110_BO6),
.D(CLBLM_R_X41Y107_SLICE_X67Y107_CO6),
.Q(CLBLM_R_X41Y107_SLICE_X67Y107_D5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf303000000000000)
  ) CLBLM_R_X41Y107_SLICE_X67Y107_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y111_SLICE_X69Y111_CO5),
.I2(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I3(CLBLM_R_X41Y110_SLICE_X67Y110_CO5),
.I4(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.I5(1'b1),
.O5(CLBLM_R_X41Y107_SLICE_X67Y107_DO5),
.O6(CLBLM_R_X41Y107_SLICE_X67Y107_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hbbfb3333bbff3333)
  ) CLBLM_R_X41Y107_SLICE_X67Y107_CLUT (
.I0(CLBLM_R_X41Y107_SLICE_X67Y107_DO6),
.I1(CLBLM_R_X41Y111_SLICE_X66Y111_BO5),
.I2(CLBLM_R_X41Y107_SLICE_X67Y107_AO6),
.I3(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.I4(CLBLM_R_X41Y107_SLICE_X67Y107_BO6),
.I5(CLBLM_R_X41Y101_SLICE_X66Y101_BO5),
.O5(CLBLM_R_X41Y107_SLICE_X67Y107_CO5),
.O6(CLBLM_R_X41Y107_SLICE_X67Y107_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000333300aa00aa)
  ) CLBLM_R_X41Y107_SLICE_X67Y107_BLUT (
.I0(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I1(CLBLL_L_X42Y103_SLICE_X69Y103_BQ),
.I2(1'b1),
.I3(CLBLM_R_X41Y107_SLICE_X66Y107_CO6),
.I4(CLBLL_L_X42Y109_SLICE_X69Y109_CO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y107_SLICE_X67Y107_BO5),
.O6(CLBLM_R_X41Y107_SLICE_X67Y107_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf070b030c0408000)
  ) CLBLM_R_X41Y107_SLICE_X67Y107_ALUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I1(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I2(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I3(CLBLM_R_X41Y107_SLICE_X66Y107_BO6),
.I4(CLBLM_R_X41Y107_SLICE_X67Y107_BO5),
.I5(CLBLM_R_X41Y106_SLICE_X66Y106_BO6),
.O5(CLBLM_R_X41Y107_SLICE_X67Y107_AO5),
.O6(CLBLM_R_X41Y107_SLICE_X67Y107_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y108_SLICE_X66Y108_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y108_SLICE_X66Y108_DO6),
.D(CLBLM_R_X41Y108_SLICE_X66Y108_CO5),
.Q(CLBLM_R_X41Y108_SLICE_X66Y108_D5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0700070000000000)
  ) CLBLM_R_X41Y108_SLICE_X66Y108_DLUT (
.I0(CLBLM_R_X41Y108_SLICE_X66Y108_CO5),
.I1(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I2(CLBLM_R_X41Y115_SLICE_X66Y115_DO6),
.I3(CLBLL_L_X42Y109_SLICE_X68Y109_DO6),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y108_SLICE_X66Y108_DO5),
.O6(CLBLM_R_X41Y108_SLICE_X66Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h080800000000c000)
  ) CLBLM_R_X41Y108_SLICE_X66Y108_CLUT (
.I0(CLBLL_L_X42Y107_SLICE_X68Y107_DO6),
.I1(CLBLM_R_X41Y108_SLICE_X67Y108_CO5),
.I2(CLBLL_L_X42Y109_SLICE_X68Y109_DQ),
.I3(CLBLL_L_X42Y109_SLICE_X68Y109_BO6),
.I4(CLBLM_R_X41Y108_SLICE_X66Y108_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X41Y108_SLICE_X66Y108_CO5),
.O6(CLBLM_R_X41Y108_SLICE_X66Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0007070700777777)
  ) CLBLM_R_X41Y108_SLICE_X66Y108_BLUT (
.I0(CLBLM_R_X41Y111_SLICE_X66Y111_AQ),
.I1(CLBLM_R_X41Y108_SLICE_X66Y108_CO5),
.I2(CLBLM_R_X41Y107_SLICE_X67Y107_D5Q),
.I3(CLBLM_R_X41Y114_SLICE_X67Y114_B5Q),
.I4(CLBLL_L_X42Y110_SLICE_X69Y110_BO5),
.I5(CLBLM_R_X41Y110_SLICE_X66Y110_DO5),
.O5(CLBLM_R_X41Y108_SLICE_X66Y108_BO5),
.O6(CLBLM_R_X41Y108_SLICE_X66Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hff02ff02fd08f500)
  ) CLBLM_R_X41Y108_SLICE_X66Y108_ALUT (
.I0(CLBLL_L_X42Y109_SLICE_X68Y109_DO6),
.I1(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I2(CLBLM_R_X41Y115_SLICE_X66Y115_DO6),
.I3(CLBLL_L_X42Y109_SLICE_X68Y109_DQ),
.I4(CLBLM_R_X41Y108_SLICE_X66Y108_CO5),
.I5(CLBLM_R_X41Y110_SLICE_X66Y110_CO6),
.O5(CLBLM_R_X41Y108_SLICE_X66Y108_AO5),
.O6(CLBLM_R_X41Y108_SLICE_X66Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y108_SLICE_X67Y108_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLM_R_X41Y108_SLICE_X67Y108_AO6),
.Q(CLBLM_R_X41Y108_SLICE_X67Y108_D5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0003000300000000)
  ) CLBLM_R_X41Y108_SLICE_X67Y108_DLUT (
.I0(1'b1),
.I1(CLBLM_R_X41Y110_SLICE_X66Y110_B5Q),
.I2(CLBLL_L_X42Y109_SLICE_X68Y109_D5Q),
.I3(CLBLL_L_X42Y102_SLICE_X68Y102_BQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y108_SLICE_X67Y108_DO5),
.O6(CLBLM_R_X41Y108_SLICE_X67Y108_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000f011111111)
  ) CLBLM_R_X41Y108_SLICE_X67Y108_CLUT (
.I0(CLBLM_R_X41Y109_SLICE_X67Y109_D5Q),
.I1(CLBLM_R_X41Y108_SLICE_X67Y108_D5Q),
.I2(CLBLL_L_X42Y108_SLICE_X68Y108_C5Q),
.I3(CLBLM_R_X41Y102_SLICE_X67Y102_C5Q),
.I4(CLBLL_L_X42Y109_SLICE_X69Y109_DQ),
.I5(1'b1),
.O5(CLBLM_R_X41Y108_SLICE_X67Y108_CO5),
.O6(CLBLM_R_X41Y108_SLICE_X67Y108_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0004000000000000)
  ) CLBLM_R_X41Y108_SLICE_X67Y108_BLUT (
.I0(CLBLM_R_X41Y109_SLICE_X66Y109_AQ),
.I1(CLBLM_R_X41Y108_SLICE_X67Y108_CO5),
.I2(CLBLM_R_X41Y108_SLICE_X66Y108_D5Q),
.I3(CLBLL_L_X42Y109_SLICE_X68Y109_DQ),
.I4(CLBLM_R_X41Y108_SLICE_X67Y108_CO6),
.I5(CLBLM_R_X41Y108_SLICE_X67Y108_DO6),
.O5(CLBLM_R_X41Y108_SLICE_X67Y108_BO5),
.O6(CLBLM_R_X41Y108_SLICE_X67Y108_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff1050efef0040)
  ) CLBLM_R_X41Y108_SLICE_X67Y108_ALUT (
.I0(CLBLM_R_X41Y115_SLICE_X66Y115_DO6),
.I1(CLBLL_L_X42Y110_SLICE_X69Y110_BO6),
.I2(CLBLL_L_X42Y109_SLICE_X68Y109_DO6),
.I3(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I4(CLBLM_R_X41Y108_SLICE_X67Y108_D5Q),
.I5(CLBLM_R_X41Y110_SLICE_X66Y110_DO5),
.O5(CLBLM_R_X41Y108_SLICE_X67Y108_AO5),
.O6(CLBLM_R_X41Y108_SLICE_X67Y108_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y109_SLICE_X66Y109_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y109_SLICE_X68Y109_DO6),
.D(CLBLM_R_X41Y109_SLICE_X66Y109_AO6),
.Q(CLBLM_R_X41Y109_SLICE_X66Y109_AQ),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000100000)
  ) CLBLM_R_X41Y109_SLICE_X66Y109_DLUT (
.I0(CLBLL_L_X42Y109_SLICE_X68Y109_DQ),
.I1(CLBLM_R_X41Y108_SLICE_X66Y108_D5Q),
.I2(CLBLM_R_X41Y108_SLICE_X67Y108_CO5),
.I3(CLBLL_L_X42Y109_SLICE_X69Y109_DQ),
.I4(CLBLM_R_X41Y109_SLICE_X66Y109_BO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y109_SLICE_X66Y109_DO5),
.O6(CLBLM_R_X41Y109_SLICE_X66Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0010000000040000)
  ) CLBLM_R_X41Y109_SLICE_X66Y109_CLUT (
.I0(CLBLL_L_X42Y102_SLICE_X68Y102_BQ),
.I1(CLBLM_R_X41Y110_SLICE_X66Y110_B5Q),
.I2(CLBLM_R_X41Y109_SLICE_X66Y109_AQ),
.I3(CLBLL_L_X42Y109_SLICE_X68Y109_D5Q),
.I4(CLBLM_R_X41Y109_SLICE_X66Y109_DO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y109_SLICE_X66Y109_CO5),
.O6(CLBLM_R_X41Y109_SLICE_X66Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h03030303aaaa0000)
  ) CLBLM_R_X41Y109_SLICE_X66Y109_BLUT (
.I0(CLBLM_R_X41Y109_SLICE_X67Y109_CO6),
.I1(CLBLL_L_X42Y108_SLICE_X68Y108_C5Q),
.I2(CLBLM_R_X41Y102_SLICE_X67Y102_C5Q),
.I3(1'b1),
.I4(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I5(1'b1),
.O5(CLBLM_R_X41Y109_SLICE_X66Y109_BO5),
.O6(CLBLM_R_X41Y109_SLICE_X66Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h33a000a000000000)
  ) CLBLM_R_X41Y109_SLICE_X66Y109_ALUT (
.I0(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I1(CLBLM_R_X41Y102_SLICE_X66Y102_BQ),
.I2(CLBLM_R_X41Y109_SLICE_X66Y109_CO6),
.I3(CLBLM_R_X41Y109_SLICE_X66Y109_CO5),
.I4(CLBLM_R_X41Y115_SLICE_X66Y115_BQ),
.I5(1'b1),
.O5(CLBLM_R_X41Y109_SLICE_X66Y109_AO5),
.O6(CLBLM_R_X41Y109_SLICE_X66Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y109_SLICE_X67Y109_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y109_SLICE_X68Y109_DO6),
.D(CLBLM_R_X41Y109_SLICE_X67Y109_DO5),
.Q(CLBLM_R_X41Y109_SLICE_X67Y109_D5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haa00aa00f8f88888)
  ) CLBLM_R_X41Y109_SLICE_X67Y109_DLUT (
.I0(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I1(CLBLM_R_X41Y110_SLICE_X66Y110_CO6),
.I2(CLBLM_R_X41Y102_SLICE_X66Y102_BQ),
.I3(CLBLM_R_X41Y104_SLICE_X66Y104_D5Q),
.I4(CLBLM_R_X41Y109_SLICE_X66Y109_CO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y109_SLICE_X67Y109_DO5),
.O6(CLBLM_R_X41Y109_SLICE_X67Y109_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h4400000000880000)
  ) CLBLM_R_X41Y109_SLICE_X67Y109_CLUT (
.I0(CLBLL_L_X42Y109_SLICE_X68Y109_DQ),
.I1(CLBLM_R_X41Y108_SLICE_X67Y108_CO5),
.I2(1'b1),
.I3(CLBLM_R_X41Y108_SLICE_X66Y108_D5Q),
.I4(CLBLL_L_X42Y109_SLICE_X68Y109_BO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y109_SLICE_X67Y109_CO5),
.O6(CLBLM_R_X41Y109_SLICE_X67Y109_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0100000000040000)
  ) CLBLM_R_X41Y109_SLICE_X67Y109_BLUT (
.I0(CLBLM_R_X41Y108_SLICE_X66Y108_D5Q),
.I1(CLBLM_R_X41Y109_SLICE_X67Y109_D5Q),
.I2(CLBLL_L_X42Y109_SLICE_X68Y109_DQ),
.I3(CLBLM_R_X41Y108_SLICE_X67Y108_D5Q),
.I4(CLBLL_L_X42Y109_SLICE_X68Y109_BO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y109_SLICE_X67Y109_BO5),
.O6(CLBLM_R_X41Y109_SLICE_X67Y109_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0015003f00000000)
  ) CLBLM_R_X41Y109_SLICE_X67Y109_ALUT (
.I0(CLBLL_L_X42Y68_SLICE_X68Y68_AQ),
.I1(CLBLL_L_X42Y110_SLICE_X68Y110_AO5),
.I2(CLBLM_R_X41Y114_SLICE_X67Y114_CQ),
.I3(CLBLM_R_X41Y109_SLICE_X67Y109_BO6),
.I4(CLBLM_R_X41Y109_SLICE_X67Y109_CO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y109_SLICE_X67Y109_AO5),
.O6(CLBLM_R_X41Y109_SLICE_X67Y109_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y110_SLICE_X66Y110_B5_FDSE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y110_SLICE_X66Y110_AO5),
.D(CLBLM_R_X41Y110_SLICE_X66Y110_BO5),
.Q(CLBLM_R_X41Y110_SLICE_X66Y110_B5Q),
.S(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000ffa0a0a0a0)
  ) CLBLM_R_X41Y110_SLICE_X66Y110_DLUT (
.I0(CLBLM_R_X41Y110_SLICE_X66Y110_CO5),
.I1(1'b1),
.I2(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I3(CLBLL_L_X42Y110_SLICE_X69Y110_BO6),
.I4(CLBLM_R_X41Y110_SLICE_X66Y110_CO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y110_SLICE_X66Y110_DO5),
.O6(CLBLM_R_X41Y110_SLICE_X66Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000002000100000)
  ) CLBLM_R_X41Y110_SLICE_X66Y110_CLUT (
.I0(CLBLM_R_X41Y109_SLICE_X67Y109_D5Q),
.I1(CLBLL_L_X42Y109_SLICE_X68Y109_DQ),
.I2(CLBLL_L_X42Y109_SLICE_X68Y109_BO6),
.I3(CLBLM_R_X41Y108_SLICE_X66Y108_D5Q),
.I4(CLBLM_R_X41Y108_SLICE_X67Y108_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X41Y110_SLICE_X66Y110_CO5),
.O6(CLBLM_R_X41Y110_SLICE_X66Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000002020)
  ) CLBLM_R_X41Y110_SLICE_X66Y110_BLUT (
.I0(CLBLM_R_X41Y110_SLICE_X66Y110_DO6),
.I1(CLBLM_R_X41Y109_SLICE_X66Y109_CO5),
.I2(CLBLL_L_X42Y109_SLICE_X69Y109_BO5),
.I3(1'b1),
.I4(CLBLM_R_X41Y109_SLICE_X66Y109_CO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y110_SLICE_X66Y110_BO5),
.O6(CLBLM_R_X41Y110_SLICE_X66Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0033003305050000)
  ) CLBLM_R_X41Y110_SLICE_X66Y110_ALUT (
.I0(CLBLM_R_X41Y115_SLICE_X66Y115_DO6),
.I1(CLBLM_R_X41Y110_SLICE_X66Y110_B5Q),
.I2(CLBLM_R_X41Y110_SLICE_X66Y110_DO5),
.I3(CLBLM_R_X41Y109_SLICE_X66Y109_AQ),
.I4(CLBLL_L_X42Y109_SLICE_X68Y109_DO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y110_SLICE_X66Y110_AO5),
.O6(CLBLM_R_X41Y110_SLICE_X66Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y110_SLICE_X67Y110_B5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y110_SLICE_X68Y110_BO6),
.D(CLBLM_R_X41Y110_SLICE_X67Y110_BO5),
.Q(CLBLM_R_X41Y110_SLICE_X67Y110_B5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000f7d5a280)
  ) CLBLM_R_X41Y110_SLICE_X67Y110_DLUT (
.I0(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I1(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I2(CLBLM_R_X41Y107_SLICE_X66Y107_BO6),
.I3(CLBLM_R_X41Y107_SLICE_X67Y107_BO5),
.I4(CLBLM_R_X41Y106_SLICE_X66Y106_BO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y110_SLICE_X67Y110_DO5),
.O6(CLBLM_R_X41Y110_SLICE_X67Y110_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000003110000)
  ) CLBLM_R_X41Y110_SLICE_X67Y110_CLUT (
.I0(CLBLL_L_X42Y101_SLICE_X69Y101_DO6),
.I1(CLBLM_R_X41Y101_SLICE_X67Y101_DQ),
.I2(CLBLL_L_X42Y106_SLICE_X68Y106_CO5),
.I3(CLBLM_R_X41Y101_SLICE_X67Y101_D5Q),
.I4(CLBLL_L_X42Y103_SLICE_X68Y103_BO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y110_SLICE_X67Y110_CO5),
.O6(CLBLM_R_X41Y110_SLICE_X67Y110_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ff20ffff)
  ) CLBLM_R_X41Y110_SLICE_X67Y110_BLUT (
.I0(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I1(CLBLL_L_X42Y110_SLICE_X68Y110_DO6),
.I2(CLBLM_R_X41Y110_SLICE_X67Y110_B5Q),
.I3(CLBLM_R_X41Y110_SLICE_X67Y110_AO6),
.I4(CLBLM_R_X41Y111_SLICE_X66Y111_CO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y110_SLICE_X67Y110_BO5),
.O6(CLBLM_R_X41Y110_SLICE_X67Y110_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000a8a8a000a8080)
  ) CLBLM_R_X41Y110_SLICE_X67Y110_ALUT (
.I0(CLBLM_R_X41Y107_SLICE_X67Y107_BO6),
.I1(CLBLM_R_X41Y110_SLICE_X67Y110_CO5),
.I2(CLBLL_L_X42Y104_SLICE_X68Y104_DQ),
.I3(CLBLL_L_X42Y111_SLICE_X69Y111_CO5),
.I4(CLBLM_R_X41Y101_SLICE_X67Y101_C5Q),
.I5(CLBLM_R_X41Y110_SLICE_X67Y110_DO5),
.O5(CLBLM_R_X41Y110_SLICE_X67Y110_AO5),
.O6(CLBLM_R_X41Y110_SLICE_X67Y110_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y111_SLICE_X66Y111_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLM_R_X41Y111_SLICE_X66Y111_AO5),
.Q(CLBLM_R_X41Y111_SLICE_X66Y111_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y111_SLICE_X66Y111_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y113_SLICE_X69Y113_D5Q),
.Q(CLBLM_R_X41Y111_SLICE_X66Y111_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y111_SLICE_X66Y111_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y113_SLICE_X69Y113_B5Q),
.Q(CLBLM_R_X41Y111_SLICE_X66Y111_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y111_SLICE_X66Y111_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLL_L_X42Y113_SLICE_X69Y113_DQ),
.Q(CLBLM_R_X41Y111_SLICE_X66Y111_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000cc000c00)
  ) CLBLM_R_X41Y111_SLICE_X66Y111_DLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y110_SLICE_X68Y110_DO6),
.I2(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I3(CLBLL_L_X42Y109_SLICE_X69Y109_BO5),
.I4(CLBLM_R_X41Y110_SLICE_X67Y110_B5Q),
.I5(1'b1),
.O5(CLBLM_R_X41Y111_SLICE_X66Y111_DO5),
.O6(CLBLM_R_X41Y111_SLICE_X66Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000070077)
  ) CLBLM_R_X41Y111_SLICE_X66Y111_CLUT (
.I0(CLBLL_L_X42Y110_SLICE_X68Y110_AO5),
.I1(CLBLM_R_X41Y115_SLICE_X67Y115_AQ),
.I2(CLBLM_R_X41Y111_SLICE_X66Y111_A5Q),
.I3(CLBLM_R_X41Y111_SLICE_X66Y111_DO5),
.I4(CLBLM_R_X41Y109_SLICE_X67Y109_CO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y111_SLICE_X66Y111_CO5),
.O6(CLBLM_R_X41Y111_SLICE_X66Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000faff0000)
  ) CLBLM_R_X41Y111_SLICE_X66Y111_BLUT (
.I0(CLBLM_R_X41Y109_SLICE_X67Y109_BO6),
.I1(1'b1),
.I2(CLBLL_L_X42Y102_SLICE_X68Y102_BO5),
.I3(CLBLL_L_X42Y109_SLICE_X69Y109_BO5),
.I4(CLBLM_R_X41Y108_SLICE_X66Y108_BO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y111_SLICE_X66Y111_BO5),
.O6(CLBLM_R_X41Y111_SLICE_X66Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ffff0000)
  ) CLBLM_R_X41Y111_SLICE_X66Y111_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X42Y113_SLICE_X69Y113_BQ),
.I5(1'b1),
.O5(CLBLM_R_X41Y111_SLICE_X66Y111_AO5),
.O6(CLBLM_R_X41Y111_SLICE_X66Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(0),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y111_SLICE_X67Y111_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLL_L_X42Y110_SLICE_X68Y110_BO6),
.D(CLBLM_R_X41Y111_SLICE_X67Y111_AO5),
.Q(CLBLM_R_X41Y111_SLICE_X67Y111_A5Q),
.R(CLBLL_L_X42Y96_SLICE_X69Y96_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000007f500000)
  ) CLBLM_R_X41Y111_SLICE_X67Y111_DLUT (
.I0(CLBLM_R_X41Y105_SLICE_X66Y105_DQ),
.I1(CLBLL_L_X42Y109_SLICE_X69Y109_BO5),
.I2(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I3(CLBLM_R_X41Y110_SLICE_X66Y110_DO6),
.I4(CLBLM_R_X41Y111_SLICE_X67Y111_CO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y111_SLICE_X67Y111_DO5),
.O6(CLBLM_R_X41Y111_SLICE_X67Y111_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000113355ff)
  ) CLBLM_R_X41Y111_SLICE_X67Y111_CLUT (
.I0(CLBLM_R_X41Y108_SLICE_X66Y108_CO5),
.I1(CLBLM_R_X41Y106_SLICE_X67Y106_AQ),
.I2(1'b1),
.I3(CLBLL_L_X42Y102_SLICE_X69Y102_AQ),
.I4(CLBLL_L_X42Y110_SLICE_X69Y110_BO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y111_SLICE_X67Y111_CO5),
.O6(CLBLM_R_X41Y111_SLICE_X67Y111_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000153f153f)
  ) CLBLM_R_X41Y111_SLICE_X67Y111_BLUT (
.I0(CLBLM_R_X41Y108_SLICE_X66Y108_CO5),
.I1(CLBLM_R_X41Y115_SLICE_X67Y115_BQ),
.I2(CLBLL_L_X42Y110_SLICE_X69Y110_BO5),
.I3(CLBLL_L_X42Y102_SLICE_X69Y102_CQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y111_SLICE_X67Y111_BO5),
.O6(CLBLM_R_X41Y111_SLICE_X67Y111_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000000ecccffff)
  ) CLBLM_R_X41Y111_SLICE_X67Y111_ALUT (
.I0(CLBLL_L_X42Y109_SLICE_X69Y109_BO5),
.I1(CLBLL_L_X42Y105_SLICE_X68Y105_AO6),
.I2(CLBLL_L_X42Y110_SLICE_X69Y110_BQ),
.I3(CLBLM_R_X41Y111_SLICE_X67Y111_A5Q),
.I4(CLBLM_R_X41Y111_SLICE_X67Y111_BO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y111_SLICE_X67Y111_AO5),
.O6(CLBLM_R_X41Y111_SLICE_X67Y111_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y114_SLICE_X66Y114_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLM_R_X41Y114_SLICE_X66Y114_BO6),
.Q(CLBLM_R_X41Y114_SLICE_X66Y114_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y114_SLICE_X66Y114_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLM_R_X41Y114_SLICE_X66Y114_CO5),
.Q(CLBLM_R_X41Y114_SLICE_X66Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y114_SLICE_X66Y114_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLM_R_X41Y114_SLICE_X66Y114_DO5),
.Q(CLBLM_R_X41Y114_SLICE_X66Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h30300000aaaaaaaa)
  ) CLBLM_R_X41Y114_SLICE_X66Y114_DLUT (
.I0(CLBLM_R_X41Y114_SLICE_X66Y114_AO6),
.I1(CLBLM_R_X41Y102_SLICE_X66Y102_BQ),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(1'b1),
.I4(CLBLL_L_X42Y97_SLICE_X69Y97_C5Q),
.I5(1'b1),
.O5(CLBLM_R_X41Y114_SLICE_X66Y114_DO5),
.O6(CLBLM_R_X41Y114_SLICE_X66Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000000f080)
  ) CLBLM_R_X41Y114_SLICE_X66Y114_CLUT (
.I0(CLBLL_L_X42Y97_SLICE_X69Y97_C5Q),
.I1(CLBLM_R_X41Y115_SLICE_X67Y115_D_XOR),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(CLBLM_R_X41Y114_SLICE_X66Y114_CQ),
.I4(CLBLM_R_X41Y115_SLICE_X66Y115_BO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y114_SLICE_X66Y114_CO5),
.O6(CLBLM_R_X41Y114_SLICE_X66Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5040104033333333)
  ) CLBLM_R_X41Y114_SLICE_X66Y114_BLUT (
.I0(CLBLM_R_X41Y115_SLICE_X66Y115_BO5),
.I1(CLBLM_R_X41Y114_SLICE_X66Y114_D5Q),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(CLBLL_L_X42Y97_SLICE_X69Y97_C5Q),
.I4(CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR),
.I5(1'b1),
.O5(CLBLM_R_X41Y114_SLICE_X66Y114_BO5),
.O6(CLBLM_R_X41Y114_SLICE_X66Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a0a0a02080808)
  ) CLBLM_R_X41Y114_SLICE_X66Y114_ALUT (
.I0(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I1(CLBLM_R_X41Y114_SLICE_X66Y114_DQ),
.I2(CLBLM_R_X41Y115_SLICE_X66Y115_BO5),
.I3(CLBLL_L_X42Y97_SLICE_X69Y97_C5Q),
.I4(CLBLM_R_X41Y114_SLICE_X66Y114_D5Q),
.I5(CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR),
.O5(CLBLM_R_X41Y114_SLICE_X66Y114_AO5),
.O6(CLBLM_R_X41Y114_SLICE_X66Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y114_SLICE_X67Y114_A5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y114_SLICE_X67Y114_AO5),
.Q(CLBLM_R_X41Y114_SLICE_X67Y114_A5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "B5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y114_SLICE_X67Y114_B5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y114_SLICE_X67Y114_BO5),
.Q(CLBLM_R_X41Y114_SLICE_X67Y114_B5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y114_SLICE_X67Y114_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y114_SLICE_X67Y114_CO5),
.Q(CLBLM_R_X41Y114_SLICE_X67Y114_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y114_SLICE_X67Y114_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y114_SLICE_X67Y114_DO5),
.Q(CLBLM_R_X41Y114_SLICE_X67Y114_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X41Y114_SLICE_X67Y114_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X41Y114_SLICE_X67Y114_D_CY, CLBLM_R_X41Y114_SLICE_X67Y114_C_CY, CLBLM_R_X41Y114_SLICE_X67Y114_B_CY, CLBLM_R_X41Y114_SLICE_X67Y114_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({CLBLM_R_X41Y114_SLICE_X67Y114_D_XOR, CLBLM_R_X41Y114_SLICE_X67Y114_C_XOR, CLBLM_R_X41Y114_SLICE_X67Y114_B_XOR, CLBLM_R_X41Y114_SLICE_X67Y114_A_XOR}),
.S({CLBLM_R_X41Y114_SLICE_X67Y114_DO6, CLBLM_R_X41Y114_SLICE_X67Y114_CO6, CLBLM_R_X41Y114_SLICE_X67Y114_BO6, CLBLM_R_X41Y114_SLICE_X67Y114_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X41Y114_SLICE_X67Y114_DLUT (
.I0(CLBLM_R_X41Y93_SLICE_X67Y93_C5Q),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X41Y116_SLICE_X66Y116_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X41Y114_SLICE_X67Y114_DO5),
.O6(CLBLM_R_X41Y114_SLICE_X67Y114_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaaaaaaa)
  ) CLBLM_R_X41Y114_SLICE_X67Y114_CLUT (
.I0(CLBLM_R_X41Y114_SLICE_X66Y114_DQ),
.I1(1'b1),
.I2(CLBLM_R_X41Y116_SLICE_X66Y116_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y114_SLICE_X67Y114_CO5),
.O6(CLBLM_R_X41Y114_SLICE_X67Y114_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0f0f0f0)
  ) CLBLM_R_X41Y114_SLICE_X67Y114_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X41Y114_SLICE_X66Y114_DQ),
.I2(CLBLM_R_X41Y116_SLICE_X66Y116_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y114_SLICE_X67Y114_BO5),
.O6(CLBLM_R_X41Y114_SLICE_X67Y114_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ffff0000)
  ) CLBLM_R_X41Y114_SLICE_X67Y114_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X41Y114_SLICE_X66Y114_BO5),
.I3(1'b1),
.I4(CLBLM_R_X41Y116_SLICE_X66Y116_D5Q),
.I5(1'b1),
.O5(CLBLM_R_X41Y114_SLICE_X67Y114_AO5),
.O6(CLBLM_R_X41Y114_SLICE_X67Y114_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y115_SLICE_X66Y115_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLM_R_X41Y115_SLICE_X66Y115_CO6),
.Q(CLBLM_R_X41Y115_SLICE_X66Y115_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y115_SLICE_X66Y115_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLM_R_X41Y115_SLICE_X66Y115_BO6),
.Q(CLBLM_R_X41Y115_SLICE_X66Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y115_SLICE_X66Y115_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLM_R_X41Y115_SLICE_X66Y115_DO5),
.Q(CLBLM_R_X41Y115_SLICE_X66Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h00002222f0f0f0f0)
  ) CLBLM_R_X41Y115_SLICE_X66Y115_DLUT (
.I0(CLBLM_R_X41Y109_SLICE_X66Y109_CO5),
.I1(CLBLM_R_X41Y115_SLICE_X66Y115_BQ),
.I2(CLBLM_R_X41Y115_SLICE_X66Y115_AO6),
.I3(1'b1),
.I4(CLBLM_R_X41Y102_SLICE_X66Y102_BQ),
.I5(1'b1),
.O5(CLBLM_R_X41Y115_SLICE_X66Y115_DO5),
.O6(CLBLM_R_X41Y115_SLICE_X66Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5400540054001000)
  ) CLBLM_R_X41Y115_SLICE_X66Y115_CLUT (
.I0(CLBLM_R_X41Y115_SLICE_X66Y115_BO5),
.I1(CLBLL_L_X42Y97_SLICE_X69Y97_C5Q),
.I2(CLBLM_R_X41Y115_SLICE_X66Y115_D5Q),
.I3(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I4(CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR),
.I5(CLBLM_R_X41Y115_SLICE_X67Y115_C_XOR),
.O5(CLBLM_R_X41Y115_SLICE_X66Y115_CO5),
.O6(CLBLM_R_X41Y115_SLICE_X66Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h30f020a055550000)
  ) CLBLM_R_X41Y115_SLICE_X66Y115_BLUT (
.I0(CLBLM_R_X41Y115_SLICE_X66Y115_BQ),
.I1(CLBLM_R_X41Y107_SLICE_X66Y107_AO6),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(CLBLL_L_X42Y103_SLICE_X68Y103_CO6),
.I4(CLBLL_L_X42Y90_SLICE_X69Y90_CQ),
.I5(1'b1),
.O5(CLBLM_R_X41Y115_SLICE_X66Y115_BO5),
.O6(CLBLM_R_X41Y115_SLICE_X66Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050404050004040)
  ) CLBLM_R_X41Y115_SLICE_X66Y115_ALUT (
.I0(CLBLM_R_X41Y115_SLICE_X66Y115_BO5),
.I1(CLBLM_R_X41Y115_SLICE_X66Y115_DQ),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR),
.I4(CLBLL_L_X42Y97_SLICE_X69Y97_C5Q),
.I5(CLBLM_R_X41Y115_SLICE_X67Y115_A_XOR),
.O5(CLBLM_R_X41Y115_SLICE_X66Y115_AO5),
.O6(CLBLM_R_X41Y115_SLICE_X66Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y115_SLICE_X67Y115_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y115_SLICE_X67Y115_AO5),
.Q(CLBLM_R_X41Y115_SLICE_X67Y115_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y115_SLICE_X67Y115_B_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y115_SLICE_X67Y115_BO5),
.Q(CLBLM_R_X41Y115_SLICE_X67Y115_BQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y115_SLICE_X67Y115_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y115_SLICE_X67Y115_CO5),
.Q(CLBLM_R_X41Y115_SLICE_X67Y115_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y115_SLICE_X67Y115_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y116_SLICE_X66Y116_DO6),
.D(CLBLM_R_X41Y115_SLICE_X67Y115_DO5),
.Q(CLBLM_R_X41Y115_SLICE_X67Y115_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X41Y115_SLICE_X67Y115_CARRY4 (
.CI(CLBLM_R_X41Y114_SLICE_X67Y114_COUT),
.CO({CLBLM_R_X41Y115_SLICE_X67Y115_COUT, CLBLM_R_X41Y115_SLICE_X67Y115_C_CY, CLBLM_R_X41Y115_SLICE_X67Y115_B_CY, CLBLM_R_X41Y115_SLICE_X67Y115_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X41Y115_SLICE_X67Y115_D_XOR, CLBLM_R_X41Y115_SLICE_X67Y115_C_XOR, CLBLM_R_X41Y115_SLICE_X67Y115_B_XOR, CLBLM_R_X41Y115_SLICE_X67Y115_A_XOR}),
.S({CLBLM_R_X41Y115_SLICE_X67Y115_DO6, CLBLM_R_X41Y115_SLICE_X67Y115_CO6, CLBLM_R_X41Y115_SLICE_X67Y115_BO6, CLBLM_R_X41Y115_SLICE_X67Y115_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacccccccc)
  ) CLBLM_R_X41Y115_SLICE_X67Y115_DLUT (
.I0(CLBLM_R_X41Y114_SLICE_X66Y114_CQ),
.I1(CLBLM_R_X41Y116_SLICE_X66Y116_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y115_SLICE_X67Y115_DO5),
.O6(CLBLM_R_X41Y115_SLICE_X67Y115_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0aaaaaaaa)
  ) CLBLM_R_X41Y115_SLICE_X67Y115_CLUT (
.I0(CLBLM_R_X41Y115_SLICE_X66Y115_DQ),
.I1(1'b1),
.I2(CLBLM_R_X41Y115_SLICE_X66Y115_D5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y115_SLICE_X67Y115_CO5),
.O6(CLBLM_R_X41Y115_SLICE_X67Y115_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0f0f0f0)
  ) CLBLM_R_X41Y115_SLICE_X67Y115_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X41Y114_SLICE_X66Y114_CQ),
.I3(1'b1),
.I4(CLBLM_R_X41Y116_SLICE_X66Y116_DQ),
.I5(1'b1),
.O5(CLBLM_R_X41Y115_SLICE_X67Y115_BO5),
.O6(CLBLM_R_X41Y115_SLICE_X67Y115_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacccccccc)
  ) CLBLM_R_X41Y115_SLICE_X67Y115_ALUT (
.I0(CLBLM_R_X41Y115_SLICE_X66Y115_DQ),
.I1(CLBLM_R_X41Y115_SLICE_X66Y115_D5Q),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y115_SLICE_X67Y115_AO5),
.O6(CLBLM_R_X41Y115_SLICE_X67Y115_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y116_SLICE_X66Y116_D5_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLM_R_X41Y116_SLICE_X66Y116_BO6),
.Q(CLBLM_R_X41Y116_SLICE_X66Y116_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y116_SLICE_X66Y116_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLM_R_X41Y116_SLICE_X66Y116_CO6),
.Q(CLBLM_R_X41Y116_SLICE_X66Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y116_SLICE_X66Y116_D_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(1'b1),
.D(CLBLM_R_X41Y116_SLICE_X66Y116_DO5),
.Q(CLBLM_R_X41Y116_SLICE_X66Y116_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hf000f000ffff0000)
  ) CLBLM_R_X41Y116_SLICE_X66Y116_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(CLBLM_R_X41Y115_SLICE_X66Y115_BO5),
.I4(CLBLM_R_X41Y116_SLICE_X66Y116_AO6),
.I5(1'b1),
.O5(CLBLM_R_X41Y116_SLICE_X66Y116_DO5),
.O6(CLBLM_R_X41Y116_SLICE_X66Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h3030202030002020)
  ) CLBLM_R_X41Y116_SLICE_X66Y116_CLUT (
.I0(CLBLM_R_X41Y116_SLICE_X66Y116_CQ),
.I1(CLBLM_R_X41Y115_SLICE_X66Y115_BO5),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(CLBLM_R_X41Y114_SLICE_X67Y114_C_XOR),
.I4(CLBLL_L_X42Y97_SLICE_X69Y97_C5Q),
.I5(CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR),
.O5(CLBLM_R_X41Y116_SLICE_X66Y116_CO5),
.O6(CLBLM_R_X41Y116_SLICE_X66Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0a0a08080a000808)
  ) CLBLM_R_X41Y116_SLICE_X66Y116_BLUT (
.I0(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I1(CLBLM_R_X41Y116_SLICE_X66Y116_D5Q),
.I2(CLBLM_R_X41Y115_SLICE_X66Y115_BO5),
.I3(CLBLM_R_X41Y114_SLICE_X67Y114_D_XOR),
.I4(CLBLL_L_X42Y97_SLICE_X69Y97_C5Q),
.I5(CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR),
.O5(CLBLM_R_X41Y116_SLICE_X66Y116_BO5),
.O6(CLBLM_R_X41Y116_SLICE_X66Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5050500040504000)
  ) CLBLM_R_X41Y116_SLICE_X66Y116_ALUT (
.I0(CLBLM_R_X41Y115_SLICE_X66Y115_BO5),
.I1(CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR),
.I2(CLBLL_L_X42Y94_SLICE_X69Y94_CQ),
.I3(CLBLL_L_X42Y97_SLICE_X69Y97_C5Q),
.I4(CLBLM_R_X41Y116_SLICE_X66Y116_DQ),
.I5(CLBLM_R_X41Y115_SLICE_X67Y115_B_XOR),
.O5(CLBLM_R_X41Y116_SLICE_X66Y116_AO5),
.O6(CLBLM_R_X41Y116_SLICE_X66Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y116_SLICE_X67Y116_A_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLM_R_X41Y116_SLICE_X67Y116_AO5),
.Q(CLBLM_R_X41Y116_SLICE_X67Y116_AQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X41Y116_SLICE_X67Y116_C_FDRE (
.C(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O),
.CE(CLBLM_R_X41Y114_SLICE_X66Y114_DO6),
.D(CLBLM_R_X41Y116_SLICE_X67Y116_CO5),
.Q(CLBLM_R_X41Y116_SLICE_X67Y116_CQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X41Y116_SLICE_X67Y116_CARRY4 (
.CI(CLBLM_R_X41Y115_SLICE_X67Y115_COUT),
.CO({CLBLM_R_X41Y116_SLICE_X67Y116_COUT, CLBLM_R_X41Y116_SLICE_X67Y116_C_CY, CLBLM_R_X41Y116_SLICE_X67Y116_B_CY, CLBLM_R_X41Y116_SLICE_X67Y116_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X41Y116_SLICE_X67Y116_D_XOR, CLBLM_R_X41Y116_SLICE_X67Y116_C_XOR, CLBLM_R_X41Y116_SLICE_X67Y116_B_XOR, CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR}),
.S({CLBLM_R_X41Y116_SLICE_X67Y116_DO6, CLBLM_R_X41Y116_SLICE_X67Y116_CO6, CLBLM_R_X41Y116_SLICE_X67Y116_BO6, CLBLM_R_X41Y116_SLICE_X67Y116_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff0007077777)
  ) CLBLM_R_X41Y116_SLICE_X67Y116_DLUT (
.I0(CLBLM_R_X41Y109_SLICE_X67Y109_CO5),
.I1(CLBLM_R_X41Y116_SLICE_X67Y116_CQ),
.I2(CLBLM_R_X41Y115_SLICE_X67Y115_CQ),
.I3(1'b0),
.I4(CLBLL_L_X42Y110_SLICE_X68Y110_AO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y116_SLICE_X67Y116_DO5),
.O6(CLBLM_R_X41Y116_SLICE_X67Y116_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00cccccccc)
  ) CLBLM_R_X41Y116_SLICE_X67Y116_CLUT (
.I0(1'b1),
.I1(CLBLL_L_X42Y113_SLICE_X69Y113_C5Q),
.I2(1'b1),
.I3(1'b0),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X41Y116_SLICE_X67Y116_CO5),
.O6(CLBLM_R_X41Y116_SLICE_X67Y116_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0113355ff)
  ) CLBLM_R_X41Y116_SLICE_X67Y116_BLUT (
.I0(CLBLM_R_X41Y109_SLICE_X67Y109_CO5),
.I1(CLBLM_R_X41Y115_SLICE_X67Y115_DQ),
.I2(1'b0),
.I3(CLBLM_R_X41Y116_SLICE_X67Y116_AQ),
.I4(CLBLL_L_X42Y110_SLICE_X68Y110_AO5),
.I5(1'b1),
.O5(CLBLM_R_X41Y116_SLICE_X67Y116_BO5),
.O6(CLBLM_R_X41Y116_SLICE_X67Y116_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaaffff0000)
  ) CLBLM_R_X41Y116_SLICE_X67Y116_ALUT (
.I0(1'b0),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLL_L_X42Y113_SLICE_X69Y113_AQ),
.I5(1'b1),
.O5(CLBLM_R_X41Y116_SLICE_X67Y116_AO5),
.O6(CLBLM_R_X41Y116_SLICE_X67Y116_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X57Y125_IOB_X1Y126_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_O),
.O(CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_O),
.O(CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_O),
.O(CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y55_IOB_X0Y55_OBUF (
.I(CLBLM_R_X3Y59_SLICE_X3Y59_B5Q),
.O(led[1])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y57_IOB_X0Y57_OBUF (
.I(CLBLM_R_X3Y60_SLICE_X3Y60_BQ),
.O(led[3])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y59_IOB_X0Y59_OBUF (
.I(CLBLM_R_X3Y60_SLICE_X3Y60_B5Q),
.O(led[2])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y67_IOB_X0Y68_OBUF (
.I(CLBLM_R_X3Y59_SLICE_X3Y59_AQ),
.O(led[0])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X57Y125_IOB_X1Y126_IBUF (
.I(clk),
.O(RIOB33_X57Y125_IOB_X1Y126_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X57Y127_IOB_X1Y127_OBUF (
.I(CLBLL_L_X42Y101_SLICE_X68Y101_A5Q),
.O(tx)
  );
  assign CLBLL_L_X42Y43_SLICE_X68Y43_A = CLBLL_L_X42Y43_SLICE_X68Y43_AO6;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_B = CLBLL_L_X42Y43_SLICE_X68Y43_BO6;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_C = CLBLL_L_X42Y43_SLICE_X68Y43_CO6;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_D = CLBLL_L_X42Y43_SLICE_X68Y43_DO6;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_BMUX = CLBLL_L_X42Y43_SLICE_X68Y43_B_XOR;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_CMUX = CLBLL_L_X42Y43_SLICE_X68Y43_C_XOR;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_DMUX = CLBLL_L_X42Y43_SLICE_X68Y43_D_XOR;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_A = CLBLL_L_X42Y43_SLICE_X69Y43_AO6;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_B = CLBLL_L_X42Y43_SLICE_X69Y43_BO6;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_C = CLBLL_L_X42Y43_SLICE_X69Y43_CO6;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_D = CLBLL_L_X42Y43_SLICE_X69Y43_DO6;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_A = CLBLL_L_X42Y68_SLICE_X68Y68_AO6;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_B = CLBLL_L_X42Y68_SLICE_X68Y68_BO6;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_C = CLBLL_L_X42Y68_SLICE_X68Y68_CO6;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_D = CLBLL_L_X42Y68_SLICE_X68Y68_DO6;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_AMUX = CLBLL_L_X42Y68_SLICE_X68Y68_A5Q;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_BMUX = CLBLL_L_X42Y68_SLICE_X68Y68_B5Q;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_CMUX = CLBLL_L_X42Y68_SLICE_X68Y68_C5Q;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_DMUX = CLBLL_L_X42Y68_SLICE_X68Y68_D5Q;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_A = CLBLL_L_X42Y68_SLICE_X69Y68_AO6;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_B = CLBLL_L_X42Y68_SLICE_X69Y68_BO6;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_C = CLBLL_L_X42Y68_SLICE_X69Y68_CO6;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_D = CLBLL_L_X42Y68_SLICE_X69Y68_DO6;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_A = CLBLL_L_X42Y69_SLICE_X68Y69_AO6;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_B = CLBLL_L_X42Y69_SLICE_X68Y69_BO6;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_C = CLBLL_L_X42Y69_SLICE_X68Y69_CO6;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_D = CLBLL_L_X42Y69_SLICE_X68Y69_DO6;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_AMUX = CLBLL_L_X42Y69_SLICE_X68Y69_AO5;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_BMUX = CLBLL_L_X42Y69_SLICE_X68Y69_B_XOR;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_CMUX = CLBLL_L_X42Y69_SLICE_X68Y69_C_XOR;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_DMUX = CLBLL_L_X42Y69_SLICE_X68Y69_D_XOR;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_A = CLBLL_L_X42Y69_SLICE_X69Y69_AO6;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_B = CLBLL_L_X42Y69_SLICE_X69Y69_BO6;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_C = CLBLL_L_X42Y69_SLICE_X69Y69_CO6;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_D = CLBLL_L_X42Y69_SLICE_X69Y69_DO6;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_CMUX = CLBLL_L_X42Y69_SLICE_X69Y69_CO5;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_A = CLBLL_L_X42Y70_SLICE_X68Y70_AO6;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_B = CLBLL_L_X42Y70_SLICE_X68Y70_BO6;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_C = CLBLL_L_X42Y70_SLICE_X68Y70_CO6;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_D = CLBLL_L_X42Y70_SLICE_X68Y70_DO6;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_AMUX = CLBLL_L_X42Y70_SLICE_X68Y70_A_XOR;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_BMUX = CLBLL_L_X42Y70_SLICE_X68Y70_B_XOR;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_CMUX = CLBLL_L_X42Y70_SLICE_X68Y70_C_XOR;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_DMUX = CLBLL_L_X42Y70_SLICE_X68Y70_D_XOR;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_A = CLBLL_L_X42Y70_SLICE_X69Y70_AO6;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_B = CLBLL_L_X42Y70_SLICE_X69Y70_BO6;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_C = CLBLL_L_X42Y70_SLICE_X69Y70_CO6;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_D = CLBLL_L_X42Y70_SLICE_X69Y70_DO6;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_A = CLBLL_L_X42Y71_SLICE_X68Y71_AO6;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_B = CLBLL_L_X42Y71_SLICE_X68Y71_BO6;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_C = CLBLL_L_X42Y71_SLICE_X68Y71_CO6;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_D = CLBLL_L_X42Y71_SLICE_X68Y71_DO6;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_AMUX = CLBLL_L_X42Y71_SLICE_X68Y71_AO6;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_BMUX = CLBLL_L_X42Y71_SLICE_X68Y71_B5Q;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_CMUX = CLBLL_L_X42Y71_SLICE_X68Y71_CO5;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_DMUX = CLBLL_L_X42Y71_SLICE_X68Y71_DO5;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_A = CLBLL_L_X42Y71_SLICE_X69Y71_AO6;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_B = CLBLL_L_X42Y71_SLICE_X69Y71_BO6;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_C = CLBLL_L_X42Y71_SLICE_X69Y71_CO6;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_D = CLBLL_L_X42Y71_SLICE_X69Y71_DO6;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_A = CLBLL_L_X42Y80_SLICE_X68Y80_AO6;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_B = CLBLL_L_X42Y80_SLICE_X68Y80_BO6;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_C = CLBLL_L_X42Y80_SLICE_X68Y80_CO6;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_D = CLBLL_L_X42Y80_SLICE_X68Y80_DO6;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_A = CLBLL_L_X42Y80_SLICE_X69Y80_AO6;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_B = CLBLL_L_X42Y80_SLICE_X69Y80_BO6;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_C = CLBLL_L_X42Y80_SLICE_X69Y80_CO6;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_D = CLBLL_L_X42Y80_SLICE_X69Y80_DO6;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_AMUX = CLBLL_L_X42Y80_SLICE_X69Y80_A5Q;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_BMUX = CLBLL_L_X42Y80_SLICE_X69Y80_B5Q;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_CMUX = CLBLL_L_X42Y80_SLICE_X69Y80_C5Q;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_DMUX = CLBLL_L_X42Y80_SLICE_X69Y80_D5Q;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_A = CLBLL_L_X42Y90_SLICE_X68Y90_AO6;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_B = CLBLL_L_X42Y90_SLICE_X68Y90_BO6;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_C = CLBLL_L_X42Y90_SLICE_X68Y90_CO6;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_D = CLBLL_L_X42Y90_SLICE_X68Y90_DO6;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_BMUX = CLBLL_L_X42Y90_SLICE_X68Y90_B_XOR;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_CMUX = CLBLL_L_X42Y90_SLICE_X68Y90_C_XOR;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_DMUX = CLBLL_L_X42Y90_SLICE_X68Y90_D_XOR;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_A = CLBLL_L_X42Y90_SLICE_X69Y90_AO6;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_B = CLBLL_L_X42Y90_SLICE_X69Y90_BO6;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_C = CLBLL_L_X42Y90_SLICE_X69Y90_CO6;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_D = CLBLL_L_X42Y90_SLICE_X69Y90_DO6;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_AMUX = CLBLL_L_X42Y90_SLICE_X69Y90_AO5;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_BMUX = CLBLL_L_X42Y90_SLICE_X69Y90_BO5;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_CMUX = CLBLL_L_X42Y90_SLICE_X69Y90_CO6;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_DMUX = CLBLL_L_X42Y90_SLICE_X69Y90_DO6;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_A = CLBLL_L_X42Y91_SLICE_X68Y91_AO6;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_B = CLBLL_L_X42Y91_SLICE_X68Y91_BO6;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_C = CLBLL_L_X42Y91_SLICE_X68Y91_CO6;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_D = CLBLL_L_X42Y91_SLICE_X68Y91_DO6;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_AMUX = CLBLL_L_X42Y91_SLICE_X68Y91_A_XOR;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_BMUX = CLBLL_L_X42Y91_SLICE_X68Y91_B_XOR;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_CMUX = CLBLL_L_X42Y91_SLICE_X68Y91_C_XOR;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_DMUX = CLBLL_L_X42Y91_SLICE_X68Y91_D_XOR;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_A = CLBLL_L_X42Y91_SLICE_X69Y91_AO6;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_B = CLBLL_L_X42Y91_SLICE_X69Y91_BO6;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_C = CLBLL_L_X42Y91_SLICE_X69Y91_CO6;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_D = CLBLL_L_X42Y91_SLICE_X69Y91_DO6;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_AMUX = CLBLL_L_X42Y91_SLICE_X69Y91_AO5;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_DMUX = CLBLL_L_X42Y91_SLICE_X69Y91_D5Q;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_A = CLBLL_L_X42Y92_SLICE_X68Y92_AO6;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_B = CLBLL_L_X42Y92_SLICE_X68Y92_BO6;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_C = CLBLL_L_X42Y92_SLICE_X68Y92_CO6;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_D = CLBLL_L_X42Y92_SLICE_X68Y92_DO6;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_AMUX = CLBLL_L_X42Y92_SLICE_X68Y92_A_XOR;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_BMUX = CLBLL_L_X42Y92_SLICE_X68Y92_B_XOR;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_CMUX = CLBLL_L_X42Y92_SLICE_X68Y92_C_XOR;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_DMUX = CLBLL_L_X42Y92_SLICE_X68Y92_D5Q;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_A = CLBLL_L_X42Y92_SLICE_X69Y92_AO6;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_B = CLBLL_L_X42Y92_SLICE_X69Y92_BO6;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_C = CLBLL_L_X42Y92_SLICE_X69Y92_CO6;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_D = CLBLL_L_X42Y92_SLICE_X69Y92_DO6;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_AMUX = CLBLL_L_X42Y92_SLICE_X69Y92_AO6;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_BMUX = CLBLL_L_X42Y92_SLICE_X69Y92_B5Q;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_CMUX = CLBLL_L_X42Y92_SLICE_X69Y92_C5Q;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_A = CLBLL_L_X42Y93_SLICE_X68Y93_AO6;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_B = CLBLL_L_X42Y93_SLICE_X68Y93_BO6;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_C = CLBLL_L_X42Y93_SLICE_X68Y93_CO6;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_D = CLBLL_L_X42Y93_SLICE_X68Y93_DO6;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_AMUX = CLBLL_L_X42Y93_SLICE_X68Y93_A5Q;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_BMUX = CLBLL_L_X42Y93_SLICE_X68Y93_B_XOR;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_CMUX = CLBLL_L_X42Y93_SLICE_X68Y93_C_XOR;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_DMUX = CLBLL_L_X42Y93_SLICE_X68Y93_D_XOR;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_A = CLBLL_L_X42Y93_SLICE_X69Y93_AO6;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_B = CLBLL_L_X42Y93_SLICE_X69Y93_BO6;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_C = CLBLL_L_X42Y93_SLICE_X69Y93_CO6;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_D = CLBLL_L_X42Y93_SLICE_X69Y93_DO6;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_AMUX = CLBLL_L_X42Y93_SLICE_X69Y93_AO6;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_BMUX = CLBLL_L_X42Y93_SLICE_X69Y93_BO5;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_CMUX = CLBLL_L_X42Y93_SLICE_X69Y93_CO5;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_DMUX = CLBLL_L_X42Y93_SLICE_X69Y93_DO6;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_A = CLBLL_L_X42Y94_SLICE_X68Y94_AO6;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_B = CLBLL_L_X42Y94_SLICE_X68Y94_BO6;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_C = CLBLL_L_X42Y94_SLICE_X68Y94_CO6;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_D = CLBLL_L_X42Y94_SLICE_X68Y94_DO6;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_AMUX = CLBLL_L_X42Y94_SLICE_X68Y94_A_XOR;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_BMUX = CLBLL_L_X42Y94_SLICE_X68Y94_B_XOR;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_CMUX = CLBLL_L_X42Y94_SLICE_X68Y94_C_XOR;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_DMUX = CLBLL_L_X42Y94_SLICE_X68Y94_D_XOR;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_A = CLBLL_L_X42Y94_SLICE_X69Y94_AO6;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_B = CLBLL_L_X42Y94_SLICE_X69Y94_BO6;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_C = CLBLL_L_X42Y94_SLICE_X69Y94_CO6;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_D = CLBLL_L_X42Y94_SLICE_X69Y94_DO6;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_AMUX = CLBLL_L_X42Y94_SLICE_X69Y94_AO5;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_BMUX = CLBLL_L_X42Y94_SLICE_X69Y94_BO5;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_DMUX = CLBLL_L_X42Y94_SLICE_X69Y94_DO6;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_A = CLBLL_L_X42Y95_SLICE_X68Y95_AO6;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_B = CLBLL_L_X42Y95_SLICE_X68Y95_BO6;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_C = CLBLL_L_X42Y95_SLICE_X68Y95_CO6;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_D = CLBLL_L_X42Y95_SLICE_X68Y95_DO6;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_AMUX = CLBLL_L_X42Y95_SLICE_X68Y95_A_XOR;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_BMUX = CLBLL_L_X42Y95_SLICE_X68Y95_B_XOR;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_CMUX = CLBLL_L_X42Y95_SLICE_X68Y95_CO5;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_DMUX = CLBLL_L_X42Y95_SLICE_X68Y95_D5Q;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_A = CLBLL_L_X42Y95_SLICE_X69Y95_AO6;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_B = CLBLL_L_X42Y95_SLICE_X69Y95_BO6;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_C = CLBLL_L_X42Y95_SLICE_X69Y95_CO6;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_D = CLBLL_L_X42Y95_SLICE_X69Y95_DO6;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_AMUX = CLBLL_L_X42Y95_SLICE_X69Y95_A5Q;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_CMUX = CLBLL_L_X42Y95_SLICE_X69Y95_CO6;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_DMUX = CLBLL_L_X42Y95_SLICE_X69Y95_D5Q;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_A = CLBLL_L_X42Y96_SLICE_X68Y96_AO6;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_B = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_C = CLBLL_L_X42Y96_SLICE_X68Y96_CO6;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_D = CLBLL_L_X42Y96_SLICE_X68Y96_DO6;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_AMUX = CLBLL_L_X42Y96_SLICE_X68Y96_AO5;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_BMUX = CLBLL_L_X42Y96_SLICE_X68Y96_BO5;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_CMUX = CLBLL_L_X42Y96_SLICE_X68Y96_CO5;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_DMUX = CLBLL_L_X42Y96_SLICE_X68Y96_DO5;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_A = CLBLL_L_X42Y96_SLICE_X69Y96_AO6;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_B = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_C = CLBLL_L_X42Y96_SLICE_X69Y96_CO6;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_D = CLBLL_L_X42Y96_SLICE_X69Y96_DO6;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_AMUX = CLBLL_L_X42Y96_SLICE_X69Y96_AO6;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_BMUX = CLBLL_L_X42Y96_SLICE_X69Y96_B5Q;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_CMUX = CLBLL_L_X42Y96_SLICE_X69Y96_CO6;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_DMUX = CLBLL_L_X42Y96_SLICE_X69Y96_DO6;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_A = CLBLL_L_X42Y97_SLICE_X68Y97_AO6;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_B = CLBLL_L_X42Y97_SLICE_X68Y97_BO6;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_C = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_D = CLBLL_L_X42Y97_SLICE_X68Y97_DO6;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_AMUX = CLBLL_L_X42Y97_SLICE_X68Y97_AO5;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_BMUX = CLBLL_L_X42Y97_SLICE_X68Y97_BO5;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_CMUX = CLBLL_L_X42Y97_SLICE_X68Y97_CO5;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_DMUX = CLBLL_L_X42Y97_SLICE_X68Y97_DO5;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_A = CLBLL_L_X42Y97_SLICE_X69Y97_AO6;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_B = CLBLL_L_X42Y97_SLICE_X69Y97_BO6;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_C = CLBLL_L_X42Y97_SLICE_X69Y97_CO6;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_D = CLBLL_L_X42Y97_SLICE_X69Y97_DO6;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_AMUX = CLBLL_L_X42Y97_SLICE_X69Y97_AO6;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_BMUX = CLBLL_L_X42Y97_SLICE_X69Y97_BO5;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_CMUX = CLBLL_L_X42Y97_SLICE_X69Y97_C5Q;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_DMUX = CLBLL_L_X42Y97_SLICE_X69Y97_DO6;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_A = CLBLL_L_X42Y98_SLICE_X68Y98_AO6;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_B = CLBLL_L_X42Y98_SLICE_X68Y98_BO6;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_C = CLBLL_L_X42Y98_SLICE_X68Y98_CO6;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_D = CLBLL_L_X42Y98_SLICE_X68Y98_DO6;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_A = CLBLL_L_X42Y98_SLICE_X69Y98_AO6;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_B = CLBLL_L_X42Y98_SLICE_X69Y98_BO6;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_C = CLBLL_L_X42Y98_SLICE_X69Y98_CO6;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_D = CLBLL_L_X42Y98_SLICE_X69Y98_DO6;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_DMUX = CLBLL_L_X42Y98_SLICE_X69Y98_D5Q;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_A = CLBLL_L_X42Y101_SLICE_X68Y101_AO6;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_B = CLBLL_L_X42Y101_SLICE_X68Y101_BO6;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_C = CLBLL_L_X42Y101_SLICE_X68Y101_CO6;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_D = CLBLL_L_X42Y101_SLICE_X68Y101_DO6;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_AMUX = CLBLL_L_X42Y101_SLICE_X68Y101_A5Q;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_A = CLBLL_L_X42Y101_SLICE_X69Y101_AO6;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_B = CLBLL_L_X42Y101_SLICE_X69Y101_BO6;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_C = CLBLL_L_X42Y101_SLICE_X69Y101_CO6;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_D = CLBLL_L_X42Y101_SLICE_X69Y101_DO6;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_AMUX = CLBLL_L_X42Y101_SLICE_X69Y101_A5Q;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_BMUX = CLBLL_L_X42Y101_SLICE_X69Y101_BO5;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_CMUX = CLBLL_L_X42Y101_SLICE_X69Y101_C5Q;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_DMUX = CLBLL_L_X42Y101_SLICE_X69Y101_D5Q;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_A = CLBLL_L_X42Y102_SLICE_X68Y102_AO6;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_B = CLBLL_L_X42Y102_SLICE_X68Y102_BO6;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_C = CLBLL_L_X42Y102_SLICE_X68Y102_CO6;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_D = CLBLL_L_X42Y102_SLICE_X68Y102_DO6;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_AMUX = CLBLL_L_X42Y102_SLICE_X68Y102_AO5;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_BMUX = CLBLL_L_X42Y102_SLICE_X68Y102_BO5;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_CMUX = CLBLL_L_X42Y102_SLICE_X68Y102_CO5;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_DMUX = CLBLL_L_X42Y102_SLICE_X68Y102_DO5;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_A = CLBLL_L_X42Y102_SLICE_X69Y102_AO6;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_B = CLBLL_L_X42Y102_SLICE_X69Y102_BO6;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_C = CLBLL_L_X42Y102_SLICE_X69Y102_CO6;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_D = CLBLL_L_X42Y102_SLICE_X69Y102_DO6;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_AMUX = CLBLL_L_X42Y102_SLICE_X69Y102_A5Q;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_BMUX = CLBLL_L_X42Y102_SLICE_X69Y102_BO5;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_CMUX = CLBLL_L_X42Y102_SLICE_X69Y102_C5Q;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_DMUX = CLBLL_L_X42Y102_SLICE_X69Y102_D5Q;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_A = CLBLL_L_X42Y103_SLICE_X68Y103_AO6;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_B = CLBLL_L_X42Y103_SLICE_X68Y103_BO6;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_C = CLBLL_L_X42Y103_SLICE_X68Y103_CO6;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_D = CLBLL_L_X42Y103_SLICE_X68Y103_DO6;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_AMUX = CLBLL_L_X42Y103_SLICE_X68Y103_AO6;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_BMUX = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_CMUX = CLBLL_L_X42Y103_SLICE_X68Y103_CO5;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_DMUX = CLBLL_L_X42Y103_SLICE_X68Y103_DO5;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_A = CLBLL_L_X42Y103_SLICE_X69Y103_AO6;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_B = CLBLL_L_X42Y103_SLICE_X69Y103_BO6;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_C = CLBLL_L_X42Y103_SLICE_X69Y103_CO6;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_D = CLBLL_L_X42Y103_SLICE_X69Y103_DO6;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_AMUX = CLBLL_L_X42Y103_SLICE_X69Y103_AO5;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_BMUX = CLBLL_L_X42Y103_SLICE_X69Y103_B_XOR;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_CMUX = CLBLL_L_X42Y103_SLICE_X69Y103_C_XOR;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_DMUX = CLBLL_L_X42Y103_SLICE_X69Y103_D_XOR;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_A = CLBLL_L_X42Y104_SLICE_X68Y104_AO6;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_B = CLBLL_L_X42Y104_SLICE_X68Y104_BO6;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_C = CLBLL_L_X42Y104_SLICE_X68Y104_CO6;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_D = CLBLL_L_X42Y104_SLICE_X68Y104_DO6;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_AMUX = CLBLL_L_X42Y104_SLICE_X68Y104_AO6;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_BMUX = CLBLL_L_X42Y104_SLICE_X68Y104_BO6;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_CMUX = CLBLL_L_X42Y104_SLICE_X68Y104_CO6;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_DMUX = CLBLL_L_X42Y104_SLICE_X68Y104_DO5;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_A = CLBLL_L_X42Y104_SLICE_X69Y104_AO6;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_B = CLBLL_L_X42Y104_SLICE_X69Y104_BO6;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_C = CLBLL_L_X42Y104_SLICE_X69Y104_CO6;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_D = CLBLL_L_X42Y104_SLICE_X69Y104_DO6;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_AMUX = CLBLL_L_X42Y104_SLICE_X69Y104_A_XOR;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_BMUX = CLBLL_L_X42Y104_SLICE_X69Y104_BO5;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_CMUX = CLBLL_L_X42Y104_SLICE_X69Y104_CO5;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_DMUX = CLBLL_L_X42Y104_SLICE_X69Y104_DO5;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_A = CLBLL_L_X42Y105_SLICE_X68Y105_AO6;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_B = CLBLL_L_X42Y105_SLICE_X68Y105_BO6;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_C = CLBLL_L_X42Y105_SLICE_X68Y105_CO6;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_D = CLBLL_L_X42Y105_SLICE_X68Y105_DO6;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_AMUX = CLBLL_L_X42Y105_SLICE_X68Y105_AO6;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_BMUX = CLBLL_L_X42Y105_SLICE_X68Y105_BO5;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_CMUX = CLBLL_L_X42Y105_SLICE_X68Y105_CO5;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_DMUX = CLBLL_L_X42Y105_SLICE_X68Y105_DO6;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_A = CLBLL_L_X42Y105_SLICE_X69Y105_AO6;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_B = CLBLL_L_X42Y105_SLICE_X69Y105_BO6;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_C = CLBLL_L_X42Y105_SLICE_X69Y105_CO6;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_D = CLBLL_L_X42Y105_SLICE_X69Y105_DO6;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_AMUX = CLBLL_L_X42Y105_SLICE_X69Y105_A5Q;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_BMUX = CLBLL_L_X42Y105_SLICE_X69Y105_BO5;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_CMUX = CLBLL_L_X42Y105_SLICE_X69Y105_CO5;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_DMUX = CLBLL_L_X42Y105_SLICE_X69Y105_DO5;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_A = CLBLL_L_X42Y106_SLICE_X68Y106_AO6;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_B = CLBLL_L_X42Y106_SLICE_X68Y106_BO6;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_C = CLBLL_L_X42Y106_SLICE_X68Y106_CO6;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_D = CLBLL_L_X42Y106_SLICE_X68Y106_DO6;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_AMUX = CLBLL_L_X42Y106_SLICE_X68Y106_A5Q;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_BMUX = CLBLL_L_X42Y106_SLICE_X68Y106_BO5;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_CMUX = CLBLL_L_X42Y106_SLICE_X68Y106_CO5;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_DMUX = CLBLL_L_X42Y106_SLICE_X68Y106_DO5;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_A = CLBLL_L_X42Y106_SLICE_X69Y106_AO6;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_B = CLBLL_L_X42Y106_SLICE_X69Y106_BO6;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_C = CLBLL_L_X42Y106_SLICE_X69Y106_CO6;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_D = CLBLL_L_X42Y106_SLICE_X69Y106_DO6;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_AMUX = CLBLL_L_X42Y106_SLICE_X69Y106_AO6;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_BMUX = CLBLL_L_X42Y106_SLICE_X69Y106_BO5;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_CMUX = CLBLL_L_X42Y106_SLICE_X69Y106_CO5;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_DMUX = CLBLL_L_X42Y106_SLICE_X69Y106_DO5;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_A = CLBLL_L_X42Y107_SLICE_X68Y107_AO6;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_B = CLBLL_L_X42Y107_SLICE_X68Y107_BO6;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_C = CLBLL_L_X42Y107_SLICE_X68Y107_CO6;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_D = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_AMUX = CLBLL_L_X42Y107_SLICE_X68Y107_AO6;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_BMUX = CLBLL_L_X42Y107_SLICE_X68Y107_BO5;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_CMUX = CLBLL_L_X42Y107_SLICE_X68Y107_CO6;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_DMUX = CLBLL_L_X42Y107_SLICE_X68Y107_DO5;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_A = CLBLL_L_X42Y107_SLICE_X69Y107_AO6;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_B = CLBLL_L_X42Y107_SLICE_X69Y107_BO6;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_C = CLBLL_L_X42Y107_SLICE_X69Y107_CO6;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_D = CLBLL_L_X42Y107_SLICE_X69Y107_DO6;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_AMUX = CLBLL_L_X42Y107_SLICE_X69Y107_A5Q;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_BMUX = CLBLL_L_X42Y107_SLICE_X69Y107_B5Q;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_CMUX = CLBLL_L_X42Y107_SLICE_X69Y107_C5Q;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_DMUX = CLBLL_L_X42Y107_SLICE_X69Y107_D5Q;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_A = CLBLL_L_X42Y108_SLICE_X68Y108_AO6;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_B = CLBLL_L_X42Y108_SLICE_X68Y108_BO6;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_C = CLBLL_L_X42Y108_SLICE_X68Y108_CO6;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_D = CLBLL_L_X42Y108_SLICE_X68Y108_DO6;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_AMUX = CLBLL_L_X42Y108_SLICE_X68Y108_AO5;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_BMUX = CLBLL_L_X42Y108_SLICE_X68Y108_BO5;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_CMUX = CLBLL_L_X42Y108_SLICE_X68Y108_C5Q;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_DMUX = CLBLL_L_X42Y108_SLICE_X68Y108_DO5;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_A = CLBLL_L_X42Y108_SLICE_X69Y108_AO6;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_B = CLBLL_L_X42Y108_SLICE_X69Y108_BO6;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_C = CLBLL_L_X42Y108_SLICE_X69Y108_CO6;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_D = CLBLL_L_X42Y108_SLICE_X69Y108_DO6;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_AMUX = CLBLL_L_X42Y108_SLICE_X69Y108_A5Q;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_BMUX = CLBLL_L_X42Y108_SLICE_X69Y108_BO5;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_CMUX = CLBLL_L_X42Y108_SLICE_X69Y108_CO5;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_DMUX = CLBLL_L_X42Y108_SLICE_X69Y108_D5Q;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_A = CLBLL_L_X42Y109_SLICE_X68Y109_AO6;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_B = CLBLL_L_X42Y109_SLICE_X68Y109_BO6;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_C = CLBLL_L_X42Y109_SLICE_X68Y109_CO6;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_D = CLBLL_L_X42Y109_SLICE_X68Y109_DO6;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_AMUX = CLBLL_L_X42Y109_SLICE_X68Y109_AO6;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_BMUX = CLBLL_L_X42Y109_SLICE_X68Y109_BO6;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_CMUX = CLBLL_L_X42Y109_SLICE_X68Y109_CO6;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_DMUX = CLBLL_L_X42Y109_SLICE_X68Y109_D5Q;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_A = CLBLL_L_X42Y109_SLICE_X69Y109_AO6;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_B = CLBLL_L_X42Y109_SLICE_X69Y109_BO6;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_C = CLBLL_L_X42Y109_SLICE_X69Y109_CO6;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_D = CLBLL_L_X42Y109_SLICE_X69Y109_DO6;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_AMUX = CLBLL_L_X42Y109_SLICE_X69Y109_AO6;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_BMUX = CLBLL_L_X42Y109_SLICE_X69Y109_BO5;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_CMUX = CLBLL_L_X42Y109_SLICE_X69Y109_CO5;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_A = CLBLL_L_X42Y110_SLICE_X68Y110_AO6;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_B = CLBLL_L_X42Y110_SLICE_X68Y110_BO6;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_C = CLBLL_L_X42Y110_SLICE_X68Y110_CO6;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_D = CLBLL_L_X42Y110_SLICE_X68Y110_DO6;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_AMUX = CLBLL_L_X42Y110_SLICE_X68Y110_AO5;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_BMUX = CLBLL_L_X42Y110_SLICE_X68Y110_BO5;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_CMUX = CLBLL_L_X42Y110_SLICE_X68Y110_C5Q;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_DMUX = CLBLL_L_X42Y110_SLICE_X68Y110_DO5;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_A = CLBLL_L_X42Y110_SLICE_X69Y110_AO6;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_B = CLBLL_L_X42Y110_SLICE_X69Y110_BO6;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_C = CLBLL_L_X42Y110_SLICE_X69Y110_CO6;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_D = CLBLL_L_X42Y110_SLICE_X69Y110_DO6;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_AMUX = CLBLL_L_X42Y110_SLICE_X69Y110_AO5;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_BMUX = CLBLL_L_X42Y110_SLICE_X69Y110_BO5;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_CMUX = CLBLL_L_X42Y110_SLICE_X69Y110_C5Q;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_DMUX = CLBLL_L_X42Y110_SLICE_X69Y110_DO5;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_A = CLBLL_L_X42Y111_SLICE_X68Y111_AO6;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_B = CLBLL_L_X42Y111_SLICE_X68Y111_BO6;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_C = CLBLL_L_X42Y111_SLICE_X68Y111_CO6;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_D = CLBLL_L_X42Y111_SLICE_X68Y111_DO6;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_AMUX = CLBLL_L_X42Y111_SLICE_X68Y111_A5Q;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_BMUX = CLBLL_L_X42Y111_SLICE_X68Y111_B5Q;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_CMUX = CLBLL_L_X42Y111_SLICE_X68Y111_C5Q;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_DMUX = CLBLL_L_X42Y111_SLICE_X68Y111_D5Q;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_A = CLBLL_L_X42Y111_SLICE_X69Y111_AO6;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_B = CLBLL_L_X42Y111_SLICE_X69Y111_BO6;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_C = CLBLL_L_X42Y111_SLICE_X69Y111_CO6;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_D = CLBLL_L_X42Y111_SLICE_X69Y111_DO6;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_AMUX = CLBLL_L_X42Y111_SLICE_X69Y111_A5Q;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_CMUX = CLBLL_L_X42Y111_SLICE_X69Y111_CO5;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_DMUX = CLBLL_L_X42Y111_SLICE_X69Y111_D5Q;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_A = CLBLL_L_X42Y112_SLICE_X68Y112_AO6;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_B = CLBLL_L_X42Y112_SLICE_X68Y112_BO6;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_C = CLBLL_L_X42Y112_SLICE_X68Y112_CO6;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_D = CLBLL_L_X42Y112_SLICE_X68Y112_DO6;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_AMUX = CLBLL_L_X42Y112_SLICE_X68Y112_A5Q;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_BMUX = CLBLL_L_X42Y112_SLICE_X68Y112_B5Q;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_CMUX = CLBLL_L_X42Y112_SLICE_X68Y112_C5Q;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_DMUX = CLBLL_L_X42Y112_SLICE_X68Y112_D5Q;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_A = CLBLL_L_X42Y112_SLICE_X69Y112_AO6;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_B = CLBLL_L_X42Y112_SLICE_X69Y112_BO6;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_C = CLBLL_L_X42Y112_SLICE_X69Y112_CO6;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_D = CLBLL_L_X42Y112_SLICE_X69Y112_DO6;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_AMUX = CLBLL_L_X42Y112_SLICE_X69Y112_AO6;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_BMUX = CLBLL_L_X42Y112_SLICE_X69Y112_BO5;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_CMUX = CLBLL_L_X42Y112_SLICE_X69Y112_C5Q;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_DMUX = CLBLL_L_X42Y112_SLICE_X69Y112_DO5;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_A = CLBLL_L_X42Y113_SLICE_X68Y113_AO6;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_B = CLBLL_L_X42Y113_SLICE_X68Y113_BO6;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_C = CLBLL_L_X42Y113_SLICE_X68Y113_CO6;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_D = CLBLL_L_X42Y113_SLICE_X68Y113_DO6;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_DMUX = CLBLL_L_X42Y113_SLICE_X68Y113_D5Q;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_A = CLBLL_L_X42Y113_SLICE_X69Y113_AO6;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_B = CLBLL_L_X42Y113_SLICE_X69Y113_BO6;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_C = CLBLL_L_X42Y113_SLICE_X69Y113_CO6;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_D = CLBLL_L_X42Y113_SLICE_X69Y113_DO6;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_AMUX = CLBLL_L_X42Y113_SLICE_X69Y113_A5Q;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_BMUX = CLBLL_L_X42Y113_SLICE_X69Y113_B5Q;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_CMUX = CLBLL_L_X42Y113_SLICE_X69Y113_C5Q;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_DMUX = CLBLL_L_X42Y113_SLICE_X69Y113_D5Q;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_A = CLBLL_L_X42Y118_SLICE_X68Y118_AO6;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_B = CLBLL_L_X42Y118_SLICE_X68Y118_BO6;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_C = CLBLL_L_X42Y118_SLICE_X68Y118_CO6;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_D = CLBLL_L_X42Y118_SLICE_X68Y118_DO6;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_A = CLBLL_L_X42Y118_SLICE_X69Y118_AO6;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_B = CLBLL_L_X42Y118_SLICE_X69Y118_BO6;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_C = CLBLL_L_X42Y118_SLICE_X69Y118_CO6;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_D = CLBLL_L_X42Y118_SLICE_X69Y118_DO6;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_AMUX = CLBLL_L_X42Y118_SLICE_X69Y118_A5Q;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_BMUX = CLBLL_L_X42Y118_SLICE_X69Y118_B5Q;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_CMUX = CLBLL_L_X42Y118_SLICE_X69Y118_C5Q;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_DMUX = CLBLL_L_X42Y118_SLICE_X69Y118_D5Q;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_A = CLBLM_R_X3Y54_SLICE_X2Y54_AO6;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_B = CLBLM_R_X3Y54_SLICE_X2Y54_BO6;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_C = CLBLM_R_X3Y54_SLICE_X2Y54_CO6;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_D = CLBLM_R_X3Y54_SLICE_X2Y54_DO6;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_A = CLBLM_R_X3Y54_SLICE_X3Y54_AO6;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_B = CLBLM_R_X3Y54_SLICE_X3Y54_BO6;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_C = CLBLM_R_X3Y54_SLICE_X3Y54_CO6;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_D = CLBLM_R_X3Y54_SLICE_X3Y54_DO6;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_AMUX = CLBLM_R_X3Y54_SLICE_X3Y54_AO5;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_BMUX = CLBLM_R_X3Y54_SLICE_X3Y54_B5Q;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_A = CLBLM_R_X3Y55_SLICE_X2Y55_AO6;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_B = CLBLM_R_X3Y55_SLICE_X2Y55_BO6;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_C = CLBLM_R_X3Y55_SLICE_X2Y55_CO6;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_D = CLBLM_R_X3Y55_SLICE_X2Y55_DO6;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_A = CLBLM_R_X3Y55_SLICE_X3Y55_AO6;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_B = CLBLM_R_X3Y55_SLICE_X3Y55_BO6;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_C = CLBLM_R_X3Y55_SLICE_X3Y55_CO6;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_D = CLBLM_R_X3Y55_SLICE_X3Y55_DO6;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_AMUX = CLBLM_R_X3Y55_SLICE_X3Y55_A_XOR;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_BMUX = CLBLM_R_X3Y55_SLICE_X3Y55_B5Q;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_CMUX = CLBLM_R_X3Y55_SLICE_X3Y55_C_XOR;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_DMUX = CLBLM_R_X3Y55_SLICE_X3Y55_D_XOR;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_A = CLBLM_R_X3Y56_SLICE_X2Y56_AO6;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_B = CLBLM_R_X3Y56_SLICE_X2Y56_BO6;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_C = CLBLM_R_X3Y56_SLICE_X2Y56_CO6;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_D = CLBLM_R_X3Y56_SLICE_X2Y56_DO6;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_A = CLBLM_R_X3Y56_SLICE_X3Y56_AO6;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_B = CLBLM_R_X3Y56_SLICE_X3Y56_BO6;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_C = CLBLM_R_X3Y56_SLICE_X3Y56_CO6;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_D = CLBLM_R_X3Y56_SLICE_X3Y56_DO6;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_AMUX = CLBLM_R_X3Y56_SLICE_X3Y56_A_XOR;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_BMUX = CLBLM_R_X3Y56_SLICE_X3Y56_B5Q;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_CMUX = CLBLM_R_X3Y56_SLICE_X3Y56_C_XOR;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_DMUX = CLBLM_R_X3Y56_SLICE_X3Y56_D_XOR;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_A = CLBLM_R_X3Y57_SLICE_X2Y57_AO6;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_B = CLBLM_R_X3Y57_SLICE_X2Y57_BO6;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_C = CLBLM_R_X3Y57_SLICE_X2Y57_CO6;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_D = CLBLM_R_X3Y57_SLICE_X2Y57_DO6;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_A = CLBLM_R_X3Y57_SLICE_X3Y57_AO6;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_B = CLBLM_R_X3Y57_SLICE_X3Y57_BO6;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_C = CLBLM_R_X3Y57_SLICE_X3Y57_CO6;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_D = CLBLM_R_X3Y57_SLICE_X3Y57_DO6;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_AMUX = CLBLM_R_X3Y57_SLICE_X3Y57_A_XOR;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_BMUX = CLBLM_R_X3Y57_SLICE_X3Y57_B5Q;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_CMUX = CLBLM_R_X3Y57_SLICE_X3Y57_C_XOR;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_DMUX = CLBLM_R_X3Y57_SLICE_X3Y57_D_XOR;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_A = CLBLM_R_X3Y58_SLICE_X2Y58_AO6;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_B = CLBLM_R_X3Y58_SLICE_X2Y58_BO6;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_C = CLBLM_R_X3Y58_SLICE_X2Y58_CO6;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_D = CLBLM_R_X3Y58_SLICE_X2Y58_DO6;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_A = CLBLM_R_X3Y58_SLICE_X3Y58_AO6;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_B = CLBLM_R_X3Y58_SLICE_X3Y58_BO6;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_C = CLBLM_R_X3Y58_SLICE_X3Y58_CO6;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_D = CLBLM_R_X3Y58_SLICE_X3Y58_DO6;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_AMUX = CLBLM_R_X3Y58_SLICE_X3Y58_A_XOR;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_BMUX = CLBLM_R_X3Y58_SLICE_X3Y58_B5Q;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_CMUX = CLBLM_R_X3Y58_SLICE_X3Y58_C_XOR;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_DMUX = CLBLM_R_X3Y58_SLICE_X3Y58_D_XOR;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_A = CLBLM_R_X3Y59_SLICE_X2Y59_AO6;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_B = CLBLM_R_X3Y59_SLICE_X2Y59_BO6;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_C = CLBLM_R_X3Y59_SLICE_X2Y59_CO6;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_D = CLBLM_R_X3Y59_SLICE_X2Y59_DO6;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_A = CLBLM_R_X3Y59_SLICE_X3Y59_AO6;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_B = CLBLM_R_X3Y59_SLICE_X3Y59_BO6;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_C = CLBLM_R_X3Y59_SLICE_X3Y59_CO6;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_D = CLBLM_R_X3Y59_SLICE_X3Y59_DO6;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_AMUX = CLBLM_R_X3Y59_SLICE_X3Y59_A_XOR;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_BMUX = CLBLM_R_X3Y59_SLICE_X3Y59_B5Q;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_CMUX = CLBLM_R_X3Y59_SLICE_X3Y59_C_XOR;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_DMUX = CLBLM_R_X3Y59_SLICE_X3Y59_D_XOR;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_A = CLBLM_R_X3Y60_SLICE_X2Y60_AO6;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_B = CLBLM_R_X3Y60_SLICE_X2Y60_BO6;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_C = CLBLM_R_X3Y60_SLICE_X2Y60_CO6;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_D = CLBLM_R_X3Y60_SLICE_X2Y60_DO6;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_A = CLBLM_R_X3Y60_SLICE_X3Y60_AO6;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_B = CLBLM_R_X3Y60_SLICE_X3Y60_BO6;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_C = CLBLM_R_X3Y60_SLICE_X3Y60_CO6;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_D = CLBLM_R_X3Y60_SLICE_X3Y60_DO6;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_AMUX = CLBLM_R_X3Y60_SLICE_X3Y60_A_XOR;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_BMUX = CLBLM_R_X3Y60_SLICE_X3Y60_B5Q;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_A = CLBLM_R_X41Y92_SLICE_X66Y92_AO6;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_B = CLBLM_R_X41Y92_SLICE_X66Y92_BO6;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_C = CLBLM_R_X41Y92_SLICE_X66Y92_CO6;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_D = CLBLM_R_X41Y92_SLICE_X66Y92_DO6;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_A = CLBLM_R_X41Y92_SLICE_X67Y92_AO6;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_B = CLBLM_R_X41Y92_SLICE_X67Y92_BO6;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_C = CLBLM_R_X41Y92_SLICE_X67Y92_CO6;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_D = CLBLM_R_X41Y92_SLICE_X67Y92_DO6;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_AMUX = CLBLM_R_X41Y92_SLICE_X67Y92_AO5;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_BMUX = CLBLM_R_X41Y92_SLICE_X67Y92_B_XOR;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_DMUX = CLBLM_R_X41Y92_SLICE_X67Y92_D_XOR;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_A = CLBLM_R_X41Y93_SLICE_X66Y93_AO6;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_B = CLBLM_R_X41Y93_SLICE_X66Y93_BO6;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_C = CLBLM_R_X41Y93_SLICE_X66Y93_CO6;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_D = CLBLM_R_X41Y93_SLICE_X66Y93_DO6;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_A = CLBLM_R_X41Y93_SLICE_X67Y93_AO6;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_B = CLBLM_R_X41Y93_SLICE_X67Y93_BO6;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_C = CLBLM_R_X41Y93_SLICE_X67Y93_CO6;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_D = CLBLM_R_X41Y93_SLICE_X67Y93_DO6;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_AMUX = CLBLM_R_X41Y93_SLICE_X67Y93_A5Q;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_BMUX = CLBLM_R_X41Y93_SLICE_X67Y93_B5Q;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_CMUX = CLBLM_R_X41Y93_SLICE_X67Y93_C5Q;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_DMUX = CLBLM_R_X41Y93_SLICE_X67Y93_D5Q;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_A = CLBLM_R_X41Y94_SLICE_X66Y94_AO6;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_B = CLBLM_R_X41Y94_SLICE_X66Y94_BO6;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_C = CLBLM_R_X41Y94_SLICE_X66Y94_CO6;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_D = CLBLM_R_X41Y94_SLICE_X66Y94_DO6;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_A = CLBLM_R_X41Y94_SLICE_X67Y94_AO6;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_B = CLBLM_R_X41Y94_SLICE_X67Y94_BO6;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_C = CLBLM_R_X41Y94_SLICE_X67Y94_CO6;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_D = CLBLM_R_X41Y94_SLICE_X67Y94_DO6;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_AMUX = CLBLM_R_X41Y94_SLICE_X67Y94_A_XOR;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_BMUX = CLBLM_R_X41Y94_SLICE_X67Y94_B5Q;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_CMUX = CLBLM_R_X41Y94_SLICE_X67Y94_C_XOR;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_DMUX = CLBLM_R_X41Y94_SLICE_X67Y94_D_XOR;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_A = CLBLM_R_X41Y95_SLICE_X66Y95_AO6;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_B = CLBLM_R_X41Y95_SLICE_X66Y95_BO6;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_C = CLBLM_R_X41Y95_SLICE_X66Y95_CO6;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_D = CLBLM_R_X41Y95_SLICE_X66Y95_DO6;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_A = CLBLM_R_X41Y95_SLICE_X67Y95_AO6;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_B = CLBLM_R_X41Y95_SLICE_X67Y95_BO6;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_C = CLBLM_R_X41Y95_SLICE_X67Y95_CO6;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_D = CLBLM_R_X41Y95_SLICE_X67Y95_DO6;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_AMUX = CLBLM_R_X41Y95_SLICE_X67Y95_A_XOR;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_BMUX = CLBLM_R_X41Y95_SLICE_X67Y95_B_XOR;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_CMUX = CLBLM_R_X41Y95_SLICE_X67Y95_C_XOR;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_DMUX = CLBLM_R_X41Y95_SLICE_X67Y95_D_XOR;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_A = CLBLM_R_X41Y100_SLICE_X66Y100_AO6;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_B = CLBLM_R_X41Y100_SLICE_X66Y100_BO6;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_C = CLBLM_R_X41Y100_SLICE_X66Y100_CO6;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_D = CLBLM_R_X41Y100_SLICE_X66Y100_DO6;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_A = CLBLM_R_X41Y100_SLICE_X67Y100_AO6;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_B = CLBLM_R_X41Y100_SLICE_X67Y100_BO6;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_C = CLBLM_R_X41Y100_SLICE_X67Y100_CO6;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_D = CLBLM_R_X41Y100_SLICE_X67Y100_DO6;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_AMUX = CLBLM_R_X41Y100_SLICE_X67Y100_A5Q;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_BMUX = CLBLM_R_X41Y100_SLICE_X67Y100_BO5;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_CMUX = CLBLM_R_X41Y100_SLICE_X67Y100_C5Q;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_DMUX = CLBLM_R_X41Y100_SLICE_X67Y100_D5Q;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_A = CLBLM_R_X41Y101_SLICE_X66Y101_AO6;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_B = CLBLM_R_X41Y101_SLICE_X66Y101_BO6;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_C = CLBLM_R_X41Y101_SLICE_X66Y101_CO6;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_D = CLBLM_R_X41Y101_SLICE_X66Y101_DO6;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_BMUX = CLBLM_R_X41Y101_SLICE_X66Y101_BO5;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_CMUX = CLBLM_R_X41Y101_SLICE_X66Y101_CO5;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_DMUX = CLBLM_R_X41Y101_SLICE_X66Y101_DO5;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_A = CLBLM_R_X41Y101_SLICE_X67Y101_AO6;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_B = CLBLM_R_X41Y101_SLICE_X67Y101_BO6;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_C = CLBLM_R_X41Y101_SLICE_X67Y101_CO6;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_D = CLBLM_R_X41Y101_SLICE_X67Y101_DO6;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_AMUX = CLBLM_R_X41Y101_SLICE_X67Y101_AO5;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_BMUX = CLBLM_R_X41Y101_SLICE_X67Y101_BO5;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_CMUX = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_DMUX = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_A = CLBLM_R_X41Y102_SLICE_X66Y102_AO6;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_B = CLBLM_R_X41Y102_SLICE_X66Y102_BO6;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_C = CLBLM_R_X41Y102_SLICE_X66Y102_CO6;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_D = CLBLM_R_X41Y102_SLICE_X66Y102_DO6;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_AMUX = CLBLM_R_X41Y102_SLICE_X66Y102_AO5;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_BMUX = CLBLM_R_X41Y102_SLICE_X66Y102_BO5;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_CMUX = CLBLM_R_X41Y102_SLICE_X66Y102_CO5;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_DMUX = CLBLM_R_X41Y102_SLICE_X66Y102_DO5;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_A = CLBLM_R_X41Y102_SLICE_X67Y102_AO6;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_B = CLBLM_R_X41Y102_SLICE_X67Y102_BO6;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_C = CLBLM_R_X41Y102_SLICE_X67Y102_CO6;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_D = CLBLM_R_X41Y102_SLICE_X67Y102_DO6;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_AMUX = CLBLM_R_X41Y102_SLICE_X67Y102_AO5;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_BMUX = CLBLM_R_X41Y102_SLICE_X67Y102_BO5;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_CMUX = CLBLM_R_X41Y102_SLICE_X67Y102_C5Q;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_DMUX = CLBLM_R_X41Y102_SLICE_X67Y102_DO5;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_A = CLBLM_R_X41Y103_SLICE_X66Y103_AO6;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_B = CLBLM_R_X41Y103_SLICE_X66Y103_BO6;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_C = CLBLM_R_X41Y103_SLICE_X66Y103_CO6;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_D = CLBLM_R_X41Y103_SLICE_X66Y103_DO6;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_BMUX = CLBLM_R_X41Y103_SLICE_X66Y103_BO5;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_CMUX = CLBLM_R_X41Y103_SLICE_X66Y103_CO5;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_A = CLBLM_R_X41Y103_SLICE_X67Y103_AO6;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_B = CLBLM_R_X41Y103_SLICE_X67Y103_BO6;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_C = CLBLM_R_X41Y103_SLICE_X67Y103_CO6;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_D = CLBLM_R_X41Y103_SLICE_X67Y103_DO6;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_AMUX = CLBLM_R_X41Y103_SLICE_X67Y103_AO6;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_BMUX = CLBLM_R_X41Y103_SLICE_X67Y103_BO6;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_CMUX = CLBLM_R_X41Y103_SLICE_X67Y103_CO5;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_DMUX = CLBLM_R_X41Y103_SLICE_X67Y103_D5Q;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_A = CLBLM_R_X41Y104_SLICE_X66Y104_AO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_B = CLBLM_R_X41Y104_SLICE_X66Y104_BO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_C = CLBLM_R_X41Y104_SLICE_X66Y104_CO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_D = CLBLM_R_X41Y104_SLICE_X66Y104_DO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_AMUX = CLBLM_R_X41Y104_SLICE_X66Y104_AO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_BMUX = CLBLM_R_X41Y104_SLICE_X66Y104_BO5;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_CMUX = CLBLM_R_X41Y104_SLICE_X66Y104_CO5;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_DMUX = CLBLM_R_X41Y104_SLICE_X66Y104_D5Q;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_A = CLBLM_R_X41Y104_SLICE_X67Y104_AO6;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_B = CLBLM_R_X41Y104_SLICE_X67Y104_BO6;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_C = CLBLM_R_X41Y104_SLICE_X67Y104_CO6;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_D = CLBLM_R_X41Y104_SLICE_X67Y104_DO6;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_AMUX = CLBLM_R_X41Y104_SLICE_X67Y104_AO6;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_BMUX = CLBLM_R_X41Y104_SLICE_X67Y104_BO5;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_CMUX = CLBLM_R_X41Y104_SLICE_X67Y104_C5Q;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_DMUX = CLBLM_R_X41Y104_SLICE_X67Y104_DO5;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_A = CLBLM_R_X41Y105_SLICE_X66Y105_AO6;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_B = CLBLM_R_X41Y105_SLICE_X66Y105_BO6;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_C = CLBLM_R_X41Y105_SLICE_X66Y105_CO6;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_D = CLBLM_R_X41Y105_SLICE_X66Y105_DO6;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_AMUX = CLBLM_R_X41Y105_SLICE_X66Y105_AO6;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_BMUX = CLBLM_R_X41Y105_SLICE_X66Y105_BO6;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_CMUX = CLBLM_R_X41Y105_SLICE_X66Y105_CO6;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_A = CLBLM_R_X41Y105_SLICE_X67Y105_AO6;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_B = CLBLM_R_X41Y105_SLICE_X67Y105_BO6;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_C = CLBLM_R_X41Y105_SLICE_X67Y105_CO6;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_D = CLBLM_R_X41Y105_SLICE_X67Y105_DO6;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_AMUX = CLBLM_R_X41Y105_SLICE_X67Y105_AO6;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_BMUX = CLBLM_R_X41Y105_SLICE_X67Y105_BO5;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_CMUX = CLBLM_R_X41Y105_SLICE_X67Y105_CO5;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_DMUX = CLBLM_R_X41Y105_SLICE_X67Y105_DO5;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_A = CLBLM_R_X41Y106_SLICE_X66Y106_AO6;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_B = CLBLM_R_X41Y106_SLICE_X66Y106_BO6;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_C = CLBLM_R_X41Y106_SLICE_X66Y106_CO6;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_D = CLBLM_R_X41Y106_SLICE_X66Y106_DO6;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_AMUX = CLBLM_R_X41Y106_SLICE_X66Y106_AO6;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_BMUX = CLBLM_R_X41Y106_SLICE_X66Y106_BO6;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_CMUX = CLBLM_R_X41Y106_SLICE_X66Y106_CO6;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_DMUX = CLBLM_R_X41Y106_SLICE_X66Y106_DO5;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_A = CLBLM_R_X41Y106_SLICE_X67Y106_AO6;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_B = CLBLM_R_X41Y106_SLICE_X67Y106_BO6;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_C = CLBLM_R_X41Y106_SLICE_X67Y106_CO6;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_D = CLBLM_R_X41Y106_SLICE_X67Y106_DO6;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_AMUX = CLBLM_R_X41Y106_SLICE_X67Y106_A5Q;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_BMUX = CLBLM_R_X41Y106_SLICE_X67Y106_BO5;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_CMUX = CLBLM_R_X41Y106_SLICE_X67Y106_C5Q;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_DMUX = CLBLM_R_X41Y106_SLICE_X67Y106_DO5;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_A = CLBLM_R_X41Y107_SLICE_X66Y107_AO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_B = CLBLM_R_X41Y107_SLICE_X66Y107_BO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_C = CLBLM_R_X41Y107_SLICE_X66Y107_CO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_D = CLBLM_R_X41Y107_SLICE_X66Y107_DO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_AMUX = CLBLM_R_X41Y107_SLICE_X66Y107_AO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_BMUX = CLBLM_R_X41Y107_SLICE_X66Y107_BO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_CMUX = CLBLM_R_X41Y107_SLICE_X66Y107_CO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_DMUX = CLBLM_R_X41Y107_SLICE_X66Y107_DO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_A = CLBLM_R_X41Y107_SLICE_X67Y107_AO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_B = CLBLM_R_X41Y107_SLICE_X67Y107_BO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_C = CLBLM_R_X41Y107_SLICE_X67Y107_CO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_D = CLBLM_R_X41Y107_SLICE_X67Y107_DO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_AMUX = CLBLM_R_X41Y107_SLICE_X67Y107_AO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_BMUX = CLBLM_R_X41Y107_SLICE_X67Y107_BO5;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_CMUX = CLBLM_R_X41Y107_SLICE_X67Y107_CO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_DMUX = CLBLM_R_X41Y107_SLICE_X67Y107_D5Q;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_A = CLBLM_R_X41Y108_SLICE_X66Y108_AO6;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_B = CLBLM_R_X41Y108_SLICE_X66Y108_BO6;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_C = CLBLM_R_X41Y108_SLICE_X66Y108_CO6;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_D = CLBLM_R_X41Y108_SLICE_X66Y108_DO6;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_AMUX = CLBLM_R_X41Y108_SLICE_X66Y108_AO6;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_BMUX = CLBLM_R_X41Y108_SLICE_X66Y108_BO6;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_CMUX = CLBLM_R_X41Y108_SLICE_X66Y108_CO5;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_DMUX = CLBLM_R_X41Y108_SLICE_X66Y108_D5Q;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_A = CLBLM_R_X41Y108_SLICE_X67Y108_AO6;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_B = CLBLM_R_X41Y108_SLICE_X67Y108_BO6;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_C = CLBLM_R_X41Y108_SLICE_X67Y108_CO6;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_D = CLBLM_R_X41Y108_SLICE_X67Y108_DO6;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_AMUX = CLBLM_R_X41Y108_SLICE_X67Y108_AO6;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_BMUX = CLBLM_R_X41Y108_SLICE_X67Y108_BO6;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_CMUX = CLBLM_R_X41Y108_SLICE_X67Y108_CO5;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_DMUX = CLBLM_R_X41Y108_SLICE_X67Y108_D5Q;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_A = CLBLM_R_X41Y109_SLICE_X66Y109_AO6;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_B = CLBLM_R_X41Y109_SLICE_X66Y109_BO6;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_C = CLBLM_R_X41Y109_SLICE_X66Y109_CO6;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_D = CLBLM_R_X41Y109_SLICE_X66Y109_DO6;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_BMUX = CLBLM_R_X41Y109_SLICE_X66Y109_BO5;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_CMUX = CLBLM_R_X41Y109_SLICE_X66Y109_CO5;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_DMUX = CLBLM_R_X41Y109_SLICE_X66Y109_DO5;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_A = CLBLM_R_X41Y109_SLICE_X67Y109_AO6;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_B = CLBLM_R_X41Y109_SLICE_X67Y109_BO6;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_C = CLBLM_R_X41Y109_SLICE_X67Y109_CO6;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_D = CLBLM_R_X41Y109_SLICE_X67Y109_DO6;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_AMUX = CLBLM_R_X41Y109_SLICE_X67Y109_AO6;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_BMUX = CLBLM_R_X41Y109_SLICE_X67Y109_BO5;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_CMUX = CLBLM_R_X41Y109_SLICE_X67Y109_CO5;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_DMUX = CLBLM_R_X41Y109_SLICE_X67Y109_D5Q;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_A = CLBLM_R_X41Y110_SLICE_X66Y110_AO6;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_B = CLBLM_R_X41Y110_SLICE_X66Y110_BO6;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_C = CLBLM_R_X41Y110_SLICE_X66Y110_CO6;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_D = CLBLM_R_X41Y110_SLICE_X66Y110_DO6;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_AMUX = CLBLM_R_X41Y110_SLICE_X66Y110_AO5;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_BMUX = CLBLM_R_X41Y110_SLICE_X66Y110_B5Q;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_CMUX = CLBLM_R_X41Y110_SLICE_X66Y110_CO5;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_DMUX = CLBLM_R_X41Y110_SLICE_X66Y110_DO5;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_A = CLBLM_R_X41Y110_SLICE_X67Y110_AO6;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_B = CLBLM_R_X41Y110_SLICE_X67Y110_BO6;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_C = CLBLM_R_X41Y110_SLICE_X67Y110_CO6;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_D = CLBLM_R_X41Y110_SLICE_X67Y110_DO6;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_AMUX = CLBLM_R_X41Y110_SLICE_X67Y110_AO6;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_BMUX = CLBLM_R_X41Y110_SLICE_X67Y110_B5Q;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_CMUX = CLBLM_R_X41Y110_SLICE_X67Y110_CO5;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_DMUX = CLBLM_R_X41Y110_SLICE_X67Y110_DO5;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_A = CLBLM_R_X41Y111_SLICE_X66Y111_AO6;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_B = CLBLM_R_X41Y111_SLICE_X66Y111_BO6;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_C = CLBLM_R_X41Y111_SLICE_X66Y111_CO6;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_D = CLBLM_R_X41Y111_SLICE_X66Y111_DO6;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_AMUX = CLBLM_R_X41Y111_SLICE_X66Y111_A5Q;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_BMUX = CLBLM_R_X41Y111_SLICE_X66Y111_BO5;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_CMUX = CLBLM_R_X41Y111_SLICE_X66Y111_CO5;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_DMUX = CLBLM_R_X41Y111_SLICE_X66Y111_DO5;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_A = CLBLM_R_X41Y111_SLICE_X67Y111_AO6;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_B = CLBLM_R_X41Y111_SLICE_X67Y111_BO6;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_C = CLBLM_R_X41Y111_SLICE_X67Y111_CO6;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_D = CLBLM_R_X41Y111_SLICE_X67Y111_DO6;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_AMUX = CLBLM_R_X41Y111_SLICE_X67Y111_A5Q;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_BMUX = CLBLM_R_X41Y111_SLICE_X67Y111_BO5;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_CMUX = CLBLM_R_X41Y111_SLICE_X67Y111_CO5;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_DMUX = CLBLM_R_X41Y111_SLICE_X67Y111_DO5;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_A = CLBLM_R_X41Y114_SLICE_X66Y114_AO6;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_B = CLBLM_R_X41Y114_SLICE_X66Y114_BO6;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_C = CLBLM_R_X41Y114_SLICE_X66Y114_CO6;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_D = CLBLM_R_X41Y114_SLICE_X66Y114_DO6;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_AMUX = CLBLM_R_X41Y114_SLICE_X66Y114_AO6;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_BMUX = CLBLM_R_X41Y114_SLICE_X66Y114_BO5;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_DMUX = CLBLM_R_X41Y114_SLICE_X66Y114_D5Q;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_A = CLBLM_R_X41Y114_SLICE_X67Y114_AO6;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_B = CLBLM_R_X41Y114_SLICE_X67Y114_BO6;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_C = CLBLM_R_X41Y114_SLICE_X67Y114_CO6;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_D = CLBLM_R_X41Y114_SLICE_X67Y114_DO6;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_AMUX = CLBLM_R_X41Y114_SLICE_X67Y114_A5Q;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_BMUX = CLBLM_R_X41Y114_SLICE_X67Y114_B5Q;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_CMUX = CLBLM_R_X41Y114_SLICE_X67Y114_C_XOR;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_DMUX = CLBLM_R_X41Y114_SLICE_X67Y114_D_XOR;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_A = CLBLM_R_X41Y115_SLICE_X66Y115_AO6;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_B = CLBLM_R_X41Y115_SLICE_X66Y115_BO6;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_C = CLBLM_R_X41Y115_SLICE_X66Y115_CO6;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_D = CLBLM_R_X41Y115_SLICE_X66Y115_DO6;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_AMUX = CLBLM_R_X41Y115_SLICE_X66Y115_AO6;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_BMUX = CLBLM_R_X41Y115_SLICE_X66Y115_BO5;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_CMUX = CLBLM_R_X41Y115_SLICE_X66Y115_CO6;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_DMUX = CLBLM_R_X41Y115_SLICE_X66Y115_D5Q;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_A = CLBLM_R_X41Y115_SLICE_X67Y115_AO6;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_B = CLBLM_R_X41Y115_SLICE_X67Y115_BO6;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_C = CLBLM_R_X41Y115_SLICE_X67Y115_CO6;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_D = CLBLM_R_X41Y115_SLICE_X67Y115_DO6;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_AMUX = CLBLM_R_X41Y115_SLICE_X67Y115_A_XOR;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_BMUX = CLBLM_R_X41Y115_SLICE_X67Y115_B_XOR;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_CMUX = CLBLM_R_X41Y115_SLICE_X67Y115_C_XOR;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_DMUX = CLBLM_R_X41Y115_SLICE_X67Y115_D_XOR;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_A = CLBLM_R_X41Y116_SLICE_X66Y116_AO6;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_B = CLBLM_R_X41Y116_SLICE_X66Y116_BO6;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_C = CLBLM_R_X41Y116_SLICE_X66Y116_CO6;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_D = CLBLM_R_X41Y116_SLICE_X66Y116_DO6;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_AMUX = CLBLM_R_X41Y116_SLICE_X66Y116_AO6;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_BMUX = CLBLM_R_X41Y116_SLICE_X66Y116_BO6;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_DMUX = CLBLM_R_X41Y116_SLICE_X66Y116_D5Q;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_A = CLBLM_R_X41Y116_SLICE_X67Y116_AO6;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_B = CLBLM_R_X41Y116_SLICE_X67Y116_BO6;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_C = CLBLM_R_X41Y116_SLICE_X67Y116_CO6;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_D = CLBLM_R_X41Y116_SLICE_X67Y116_DO6;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_AMUX = CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_BMUX = CLBLM_R_X41Y116_SLICE_X67Y116_BO5;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_DMUX = CLBLM_R_X41Y116_SLICE_X67Y116_DO5;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_OQ = CLBLM_R_X3Y59_SLICE_X3Y59_B5Q;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_TQ = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_OQ = CLBLM_R_X3Y60_SLICE_X3Y60_B5Q;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_TQ = 1'b1;
  assign LIOI3_X0Y67_OLOGIC_X0Y68_OQ = CLBLM_R_X3Y59_SLICE_X3Y59_AQ;
  assign LIOI3_X0Y67_OLOGIC_X0Y68_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_OQ = CLBLM_R_X3Y60_SLICE_X3Y60_BQ;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_TQ = 1'b1;
  assign RIOI3_X57Y125_ILOGIC_X1Y126_O = RIOB33_X57Y125_IOB_X1Y126_I;
  assign RIOI3_X57Y127_OLOGIC_X1Y127_OQ = CLBLL_L_X42Y101_SLICE_X68Y101_A5Q;
  assign RIOI3_X57Y127_OLOGIC_X1Y127_TQ = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_A1 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_A2 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_A3 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_A4 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_A5 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_A6 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_B1 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_B2 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_B3 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_B4 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_B5 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_B6 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_C1 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_C2 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_C3 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_C4 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_C5 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_C6 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_CE = CLBLL_L_X42Y96_SLICE_X68Y96_CO5;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_D1 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_D2 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_D3 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_D4 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_D5 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_D6 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_DX = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y113_SLICE_X68Y113_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_A1 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_A2 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_A3 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_A4 = CLBLL_L_X42Y93_SLICE_X68Y93_CQ;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_A5 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_A6 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_AX = CLBLL_L_X42Y93_SLICE_X68Y93_BQ;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_B1 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_B2 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_B3 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_B4 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_B5 = CLBLL_L_X42Y93_SLICE_X68Y93_DQ;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_B6 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_BX = CLBLL_L_X42Y97_SLICE_X68Y97_AQ;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_C1 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_C2 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_C3 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_C4 = CLBLL_L_X42Y93_SLICE_X69Y93_BQ;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_C5 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_C6 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_CE = CLBLL_L_X42Y97_SLICE_X69Y97_CO6;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_CX = CLBLL_L_X42Y104_SLICE_X69Y104_CQ;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_D1 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_D2 = CLBLL_L_X42Y104_SLICE_X69Y104_AQ;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_D3 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_D4 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_D5 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_D6 = 1'b1;
  assign CLBLL_L_X42Y113_SLICE_X69Y113_DX = CLBLL_L_X42Y104_SLICE_X69Y104_BQ;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_A1 = CLBLM_R_X41Y93_SLICE_X67Y93_D5Q;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_A2 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_A3 = CLBLM_R_X41Y93_SLICE_X67Y93_A5Q;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_A4 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_A5 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_A6 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_AX = 1'b0;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_B1 = CLBLM_R_X41Y93_SLICE_X67Y93_D5Q;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_B2 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_B3 = CLBLM_R_X41Y93_SLICE_X67Y93_B5Q;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_B4 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_B5 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_B6 = 1'b1;
  assign RIOB33_X57Y127_IOB_X1Y127_O = CLBLL_L_X42Y101_SLICE_X68Y101_A5Q;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_BX = 1'b0;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_C1 = CLBLM_R_X41Y93_SLICE_X67Y93_B5Q;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_C2 = CLBLM_R_X41Y93_SLICE_X67Y93_A5Q;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_C3 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_C4 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_C5 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_C6 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_CE = CLBLM_R_X41Y116_SLICE_X66Y116_DO6;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_CIN = CLBLM_R_X41Y94_SLICE_X67Y94_COUT;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_CX = 1'b0;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_D1 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_D2 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_D3 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_D4 = CLBLM_R_X41Y93_SLICE_X67Y93_C5Q;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_D5 = CLBLM_R_X41Y94_SLICE_X67Y94_AQ;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_D6 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X67Y95_DX = 1'b0;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_A1 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_A2 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_A3 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_A4 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_A5 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_A6 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_B1 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_B2 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_B3 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_B4 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_B5 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_B6 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_C1 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_C2 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_C3 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_C4 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_C5 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_C6 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_D1 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_D2 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_D3 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_D4 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_D5 = 1'b1;
  assign CLBLM_R_X41Y95_SLICE_X66Y95_D6 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_C2 = 1'b1;
  assign CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_CE = 1'b1;
  assign CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_CE = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_C3 = CLBLM_R_X41Y116_SLICE_X66Y116_CQ;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_B3 = CLBLL_L_X42Y102_SLICE_X68Y102_CO6;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_B6 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_C1 = CLBLL_L_X42Y109_SLICE_X69Y109_CO6;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_C2 = CLBLM_R_X41Y109_SLICE_X67Y109_CO6;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_C3 = CLBLL_L_X42Y103_SLICE_X68Y103_CO6;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_C6 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_D3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_D5 = CLBLM_R_X41Y102_SLICE_X67Y102_BO5;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_D6 = 1'b1;
  assign CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_I = CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_O;
  assign CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_I = CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_O;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_C3 = CLBLM_R_X41Y115_SLICE_X66Y115_DO6;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_C4 = CLBLM_R_X41Y102_SLICE_X66Y102_CO6;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_C5 = CLBLM_R_X41Y107_SLICE_X66Y107_AO6;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_A1 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_A2 = CLBLL_L_X42Y90_SLICE_X69Y90_BO5;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_A3 = CLBLL_L_X42Y91_SLICE_X69Y91_AO5;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_A4 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_A5 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_A6 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_AX = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_B1 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_B2 = CLBLL_L_X42Y90_SLICE_X68Y90_BQ;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_B3 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_B4 = CLBLL_L_X42Y90_SLICE_X69Y90_CO6;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_B5 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_B6 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_BX = 1'b0;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_C1 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_C2 = CLBLL_L_X42Y90_SLICE_X68Y90_DQ;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_C3 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_C4 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_C5 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_C6 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_D2 = CLBLM_R_X41Y108_SLICE_X67Y108_BO6;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_CX = 1'b0;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_D1 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_D2 = CLBLL_L_X42Y90_SLICE_X69Y90_DO6;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_D3 = CLBLL_L_X42Y90_SLICE_X68Y90_AQ;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_D4 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_D5 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_D6 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X68Y90_DX = 1'b0;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_A1 = CLBLL_L_X42Y91_SLICE_X68Y91_AQ;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_A2 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_A3 = CLBLL_L_X42Y91_SLICE_X68Y91_A_XOR;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_A4 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_A5 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_A6 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_B1 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_B2 = CLBLL_L_X42Y90_SLICE_X68Y90_D_XOR;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_B3 = CLBLL_L_X42Y90_SLICE_X68Y90_AQ;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_B4 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_B5 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_B6 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_C1 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_C2 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_C3 = CLBLL_L_X42Y90_SLICE_X68Y90_BQ;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_C4 = CLBLL_L_X42Y90_SLICE_X68Y90_B_XOR;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_C5 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_C6 = 1'b1;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_CE = CLBLL_L_X42Y96_SLICE_X68Y96_AO6;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_CX = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_D1 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_D2 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_D3 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_D4 = CLBLL_L_X42Y90_SLICE_X68Y90_C_XOR;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_D5 = CLBLL_L_X42Y90_SLICE_X68Y90_DQ;
  assign CLBLL_L_X42Y90_SLICE_X69Y90_D6 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_B6 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_C2 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_D4 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_A1 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_A2 = CLBLL_L_X42Y91_SLICE_X68Y91_AQ;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_A3 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_A4 = CLBLL_L_X42Y90_SLICE_X69Y90_AO5;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_A5 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_A6 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_AX = 1'b0;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_B1 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_B2 = CLBLL_L_X42Y91_SLICE_X68Y91_BQ;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_B3 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_B4 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_B5 = CLBLL_L_X42Y94_SLICE_X69Y94_DO6;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_B6 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_BX = 1'b0;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_C1 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_C2 = CLBLL_L_X42Y91_SLICE_X68Y91_CQ;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_C3 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_C4 = CLBLL_L_X42Y94_SLICE_X69Y94_BO5;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_C5 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_C6 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_CIN = CLBLL_L_X42Y90_SLICE_X68Y90_COUT;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_CX = 1'b0;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_D1 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_D2 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_D3 = CLBLL_L_X42Y91_SLICE_X68Y91_DQ;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_D4 = CLBLL_L_X42Y94_SLICE_X69Y94_AO5;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_D5 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_D6 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X68Y91_DX = 1'b0;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_A1 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_A2 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_A3 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_A4 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_A5 = CLBLL_L_X42Y94_SLICE_X68Y94_BQ;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_A6 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_AX = CLBLL_L_X42Y91_SLICE_X69Y91_BQ;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_B1 = CLBLL_L_X42Y91_SLICE_X69Y91_BQ;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_B2 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_B3 = CLBLL_L_X42Y96_SLICE_X68Y96_AO5;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_B4 = CLBLL_L_X42Y93_SLICE_X68Y93_D_XOR;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_B5 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_B6 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_C1 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_C2 = CLBLL_L_X42Y96_SLICE_X68Y96_AO5;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_C3 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_C4 = CLBLL_L_X42Y94_SLICE_X68Y94_C_XOR;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_C5 = CLBLL_L_X42Y91_SLICE_X69Y91_CQ;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_C6 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_D1 = CLBLL_L_X42Y91_SLICE_X69Y91_DQ;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_D2 = CLBLL_L_X42Y94_SLICE_X68Y94_B_XOR;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_D3 = CLBLL_L_X42Y96_SLICE_X68Y96_AO5;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_D4 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_D5 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_D6 = 1'b1;
  assign CLBLL_L_X42Y91_SLICE_X69Y91_DX = CLBLL_L_X42Y91_SLICE_X69Y91_DQ;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_A1 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_A2 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_A3 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_A4 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_A5 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_A6 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_B1 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_B2 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_B3 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_B4 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_B5 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_B6 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_C1 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_C2 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_C3 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_C4 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_C5 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_C6 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_D1 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_D2 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_D3 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_D4 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_D5 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X68Y118_D6 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_A1 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_A2 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_A3 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_A4 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_A5 = CLBLM_R_X41Y111_SLICE_X67Y111_A5Q;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_A6 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_AX = CLBLM_R_X41Y105_SLICE_X66Y105_DQ;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_B1 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_B2 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_B3 = CLBLM_R_X41Y104_SLICE_X66Y104_D5Q;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_B4 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_B5 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_B6 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_BX = CLBLM_R_X41Y103_SLICE_X67Y103_D5Q;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_C1 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_C2 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_C3 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_C4 = CLBLM_R_X41Y107_SLICE_X67Y107_D5Q;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_C5 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_C6 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_CE = CLBLL_L_X42Y112_SLICE_X69Y112_DO5;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_CX = CLBLM_R_X41Y104_SLICE_X67Y104_C5Q;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_D1 = CLBLL_L_X42Y110_SLICE_X68Y110_C5Q;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_D2 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_D3 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_D4 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_D5 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_D6 = 1'b1;
  assign CLBLL_L_X42Y118_SLICE_X69Y118_DX = CLBLM_R_X41Y110_SLICE_X67Y110_B5Q;
  assign RIOI3_X57Y125_ILOGIC_X1Y126_D = RIOB33_X57Y125_IOB_X1Y126_I;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_A1 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_A2 = BRAM_L_X44Y95_RAMB18_X2Y38_DO12;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_A3 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_A4 = CLBLL_L_X42Y92_SLICE_X69Y92_C5Q;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_A5 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_A6 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_AX = 1'b0;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_B1 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_B2 = CLBLL_L_X42Y92_SLICE_X69Y92_AQ;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_B3 = CLBLL_L_X42Y92_SLICE_X69Y92_DQ;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_B4 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_B5 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_B6 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_BX = 1'b0;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_C1 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_C2 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_C3 = 1'b0;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_C4 = BRAM_L_X44Y95_RAMB18_X2Y38_DO14;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_C5 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_C6 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_CE = CLBLL_L_X42Y97_SLICE_X69Y97_CO6;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_CIN = CLBLL_L_X42Y91_SLICE_X68Y91_COUT;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_CX = 1'b0;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_D1 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_D2 = 1'b0;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_D3 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_D4 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_D5 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_D6 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X68Y92_DX = CLBLL_L_X42Y92_SLICE_X69Y92_C5Q;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_A1 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_A2 = CLBLM_R_X41Y93_SLICE_X67Y93_AQ;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_A3 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_A4 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_A5 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_A6 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_AX = CLBLM_R_X41Y92_SLICE_X67Y92_BQ;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_B1 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_B2 = CLBLM_R_X41Y107_SLICE_X66Y107_DO6;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_B3 = CLBLM_R_X41Y103_SLICE_X67Y103_BO6;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_B4 = CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_B5 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_B6 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_A1 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_A2 = CLBLL_L_X42Y94_SLICE_X68Y94_A_XOR;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_A3 = CLBLL_L_X42Y96_SLICE_X68Y96_AO5;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_A4 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_A5 = CLBLL_L_X42Y92_SLICE_X69Y92_BQ;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_A6 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_BX = CLBLM_R_X41Y94_SLICE_X67Y94_B5Q;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_C1 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_C2 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_B1 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_B2 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_B3 = CLBLL_L_X42Y95_SLICE_X68Y95_D5Q;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_B4 = CLBLL_L_X42Y92_SLICE_X69Y92_B5Q;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_B5 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_B6 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_C4 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_C5 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_BX = CLBLL_L_X42Y92_SLICE_X69Y92_AO6;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_CE = CLBLM_R_X41Y116_SLICE_X66Y116_DO6;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_C1 = CLBLL_L_X42Y92_SLICE_X69Y92_C5Q;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_C2 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_C3 = CLBLL_L_X42Y92_SLICE_X68Y92_A_XOR;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_C4 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_C5 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_C6 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_CX = CLBLM_R_X41Y93_SLICE_X67Y93_CQ;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_D1 = CLBLM_R_X41Y92_SLICE_X67Y92_DQ;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_D2 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_D3 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_D4 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_A1 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_A2 = 1'b1;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_D1 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_D2 = CLBLL_L_X42Y92_SLICE_X68Y92_B_XOR;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_D3 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_D4 = CLBLL_L_X42Y92_SLICE_X69Y92_DQ;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_D5 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y92_SLICE_X69Y92_D6 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_A5 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_A6 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_B1 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_B2 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_B3 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_B4 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_B5 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_B6 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_C1 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_C2 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_C3 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_C4 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_C5 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_C6 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_D1 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_D2 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_D3 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_D4 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_D5 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_D6 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_A1 = CLBLL_L_X42Y92_SLICE_X68Y92_C_XOR;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_A2 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_A3 = CLBLL_L_X42Y96_SLICE_X68Y96_BO5;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_A4 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_A5 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_A6 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_AX = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_B1 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_B2 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_B3 = CLBLL_L_X42Y97_SLICE_X68Y97_BQ;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_B4 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_B5 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_B6 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_BX = 1'b0;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_C1 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_C2 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_C3 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_C4 = CLBLL_L_X42Y95_SLICE_X69Y95_BQ;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_C5 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_C6 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_CE = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_CX = 1'b0;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_D1 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_D2 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_D3 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_D4 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_D5 = CLBLL_L_X42Y91_SLICE_X69Y91_BQ;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_D6 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_DX = 1'b0;
  assign CLBLL_L_X42Y93_SLICE_X68Y93_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_A1 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_A2 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_A3 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_A4 = CLBLL_L_X42Y110_SLICE_X68Y110_BO5;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_A5 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_A6 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_B1 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_A1 = CLBLL_L_X42Y91_SLICE_X69Y91_AQ;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_A2 = CLBLL_L_X42Y93_SLICE_X69Y93_BQ;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_A3 = BRAM_L_X44Y95_RAMB18_X2Y38_DO6;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_A4 = BRAM_L_X44Y95_RAMB18_X2Y38_DO1;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_A5 = BRAM_L_X44Y95_RAMB18_X2Y38_DO3;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_A6 = CLBLL_L_X42Y97_SLICE_X68Y97_AQ;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_B2 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_B3 = CLBLL_L_X42Y107_SLICE_X68Y107_AO6;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_B4 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_B1 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_B2 = BRAM_L_X44Y95_RAMB18_X2Y38_DO11;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_B3 = BRAM_L_X44Y95_RAMB18_X2Y38_DO14;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_B4 = BRAM_L_X44Y95_RAMB18_X2Y38_DO13;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_B5 = BRAM_L_X44Y95_RAMB18_X2Y38_DO12;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_B6 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_C1 = 1'b1;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_BX = CLBLL_L_X42Y91_SLICE_X69Y91_CQ;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_C2 = CLBLL_L_X42Y110_SLICE_X68Y110_BO5;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_C1 = CLBLL_L_X42Y96_SLICE_X68Y96_DQ;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_C2 = CLBLL_L_X42Y93_SLICE_X69Y93_AO6;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_C3 = BRAM_L_X44Y95_RAMB18_X2Y38_DO8;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_C4 = CLBLL_L_X42Y93_SLICE_X69Y93_DO6;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_C5 = CLBLL_L_X42Y95_SLICE_X68Y95_CO5;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_C6 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_CX = CLBLM_R_X41Y101_SLICE_X67Y101_AO6;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_D1 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_D2 = CLBLL_L_X42Y105_SLICE_X69Y105_DO5;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_D3 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_D4 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_D5 = CLBLM_R_X41Y101_SLICE_X67Y101_AO5;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_D1 = CLBLL_L_X42Y92_SLICE_X69Y92_AQ;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_D2 = CLBLL_L_X42Y96_SLICE_X68Y96_AQ;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_D3 = BRAM_L_X44Y95_RAMB18_X2Y38_DO4;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_D4 = CLBLL_L_X42Y93_SLICE_X69Y93_BO5;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_D5 = BRAM_L_X44Y95_RAMB18_X2Y38_DO0;
  assign CLBLL_L_X42Y93_SLICE_X69Y93_D6 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_A1 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_A2 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_A3 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_A4 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_A5 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_A6 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_B1 = CLBLM_R_X41Y105_SLICE_X67Y105_CO6;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_B2 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_B3 = CLBLL_L_X42Y107_SLICE_X68Y107_AO6;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_B4 = CLBLM_R_X41Y104_SLICE_X66Y104_DO6;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_B5 = CLBLM_R_X41Y101_SLICE_X66Y101_CO5;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_B6 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_C1 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_C2 = CLBLM_R_X41Y105_SLICE_X66Y105_CO6;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_C3 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_C4 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_C5 = CLBLM_R_X41Y105_SLICE_X67Y105_AO6;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_C6 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_D1 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_D2 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_D3 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_D4 = CLBLM_R_X41Y110_SLICE_X66Y110_DO5;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_D5 = CLBLL_L_X42Y110_SLICE_X68Y110_BO6;
  assign CLBLM_R_X41Y101_SLICE_X66Y101_D6 = 1'b1;
  assign RIOI3_X57Y127_OLOGIC_X1Y127_D1 = CLBLL_L_X42Y101_SLICE_X68Y101_A5Q;
  assign RIOI3_X57Y127_OLOGIC_X1Y127_T1 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_A2 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_A3 = CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_A1 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_A2 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_A3 = CLBLL_L_X42Y92_SLICE_X69Y92_BQ;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_A4 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_A5 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_A6 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_B3 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_B4 = CLBLL_L_X42Y105_SLICE_X69Y105_BO5;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_AX = 1'b0;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_B1 = CLBLL_L_X42Y91_SLICE_X69Y91_AO6;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_B2 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_B3 = CLBLL_L_X42Y91_SLICE_X69Y91_DQ;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_B4 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_B5 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_B6 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_B5 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_B6 = CLBLL_L_X42Y101_SLICE_X69Y101_DO6;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_BX = 1'b0;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_C1 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_C2 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_C3 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_C4 = CLBLL_L_X42Y91_SLICE_X69Y91_CQ;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_C5 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_C6 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_CIN = CLBLL_L_X42Y93_SLICE_X68Y93_COUT;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_CX = 1'b0;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_D1 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_D2 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_D3 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_D4 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_D5 = CLBLL_L_X42Y95_SLICE_X69Y95_DQ;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_D6 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X68Y94_DX = 1'b0;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_A1 = CLBLM_R_X41Y115_SLICE_X66Y115_DO6;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_A2 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_A3 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_A4 = CLBLM_R_X41Y109_SLICE_X66Y109_BO5;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_A5 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_A6 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_A1 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_A2 = CLBLL_L_X42Y91_SLICE_X68Y91_D_XOR;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_A3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_A4 = CLBLL_L_X42Y91_SLICE_X68Y91_DQ;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_A5 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_A6 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_B1 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_B2 = CLBLM_R_X41Y102_SLICE_X66Y102_BO5;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_B1 = CLBLL_L_X42Y91_SLICE_X68Y91_CQ;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_B2 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_B3 = CLBLL_L_X42Y91_SLICE_X68Y91_C_XOR;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_B4 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_B5 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_B6 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_B4 = CLBLL_L_X42Y102_SLICE_X68Y102_DO6;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_B5 = CLBLL_L_X42Y103_SLICE_X68Y103_CO6;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_C1 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_C2 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_C3 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_C4 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_C5 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_C6 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_C4 = CLBLM_R_X41Y102_SLICE_X66Y102_BO5;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_C5 = 1'b1;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_CE = CLBLM_R_X41Y102_SLICE_X67Y102_AO5;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_D1 = CLBLM_R_X41Y109_SLICE_X66Y109_BO5;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_CX = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_D2 = CLBLM_R_X41Y108_SLICE_X67Y108_BO6;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_D1 = CLBLL_L_X42Y91_SLICE_X68Y91_BQ;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_D2 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_D3 = CLBLL_L_X42Y91_SLICE_X68Y91_B_XOR;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_D4 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_D5 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y94_SLICE_X69Y94_D6 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X67Y102_D4 = CLBLL_L_X42Y109_SLICE_X69Y109_BO5;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_A1 = CLBLM_R_X41Y102_SLICE_X66Y102_CO5;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_A2 = CLBLL_L_X42Y109_SLICE_X69Y109_CO6;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_A3 = CLBLM_R_X41Y109_SLICE_X67Y109_CO6;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_A4 = CLBLM_R_X41Y102_SLICE_X66Y102_BO5;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_A5 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_A6 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_B1 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_B2 = CLBLL_L_X42Y102_SLICE_X68Y102_AO6;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_B3 = CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_B4 = CLBLM_R_X41Y105_SLICE_X67Y105_CO6;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_B5 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_B6 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_A1 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_A2 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_A3 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_A4 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_A5 = CLBLL_L_X42Y80_SLICE_X69Y80_CQ;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_A6 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_BX = CLBLM_R_X41Y102_SLICE_X66Y102_DO5;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_C1 = CLBLL_L_X42Y103_SLICE_X68Y103_CO6;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_AX = CLBLL_L_X42Y80_SLICE_X69Y80_D5Q;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_C2 = CLBLM_R_X41Y108_SLICE_X67Y108_BO6;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_B1 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_B2 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_B3 = CLBLL_L_X42Y101_SLICE_X69Y101_BQ;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_B4 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_B5 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_B6 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_C6 = 1'b1;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_BX = CLBLL_L_X42Y80_SLICE_X69Y80_C5Q;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_C1 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_C2 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_C3 = CLBLL_L_X42Y80_SLICE_X69Y80_BQ;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_C4 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_C5 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_C6 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_CE = CLBLM_R_X41Y114_SLICE_X66Y114_DO6;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_D1 = CLBLL_L_X42Y103_SLICE_X68Y103_CO6;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_D3 = CLBLL_L_X42Y97_SLICE_X69Y97_C5Q;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_D4 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_D5 = CLBLM_R_X41Y102_SLICE_X66Y102_BQ;
  assign CLBLM_R_X41Y102_SLICE_X66Y102_D6 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_CX = CLBLL_L_X42Y80_SLICE_X69Y80_DQ;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_D1 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_D2 = CLBLL_L_X42Y80_SLICE_X69Y80_A5Q;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_D3 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_D4 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_D5 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_D6 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X68Y68_DX = CLBLL_L_X42Y80_SLICE_X69Y80_AQ;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_A1 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_A2 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_A3 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_A4 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_A5 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_A6 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_B1 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_B2 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_B3 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_B4 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_B5 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_B6 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_C1 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_C2 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_C3 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_C4 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_C5 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_C6 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_D1 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_D2 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_D3 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_D4 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_D5 = 1'b1;
  assign CLBLL_L_X42Y68_SLICE_X69Y68_D6 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_C3 = CLBLM_R_X41Y104_SLICE_X67Y104_C5Q;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_A1 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_A2 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_A3 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_A4 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_A5 = CLBLL_L_X42Y95_SLICE_X69Y95_A5Q;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_A6 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_C5 = CLBLM_R_X41Y103_SLICE_X66Y103_BO5;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_C6 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_AX = 1'b0;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_B1 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_B2 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_B3 = CLBLL_L_X42Y96_SLICE_X68Y96_CQ;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_B4 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_B5 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_B6 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_BX = 1'b0;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_C1 = CLBLL_L_X42Y96_SLICE_X68Y96_AQ;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_C2 = BRAM_L_X44Y95_RAMB18_X2Y38_DO0;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_C3 = 1'b0;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_C4 = CLBLL_L_X42Y95_SLICE_X69Y95_D5Q;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_C5 = BRAM_L_X44Y95_RAMB18_X2Y38_DO7;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_C6 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_CIN = CLBLL_L_X42Y94_SLICE_X68Y94_COUT;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_CX = 1'b0;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_D1 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_D2 = 1'b0;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_D3 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_D4 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_D5 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_D6 = 1'b1;
  assign CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_CE = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X68Y95_DX = CLBLL_L_X42Y95_SLICE_X69Y95_AO6;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_A1 = CLBLM_R_X41Y107_SLICE_X67Y107_BO6;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_A1 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_A2 = 1'b1;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_A3 = CLBLL_L_X42Y95_SLICE_X68Y95_D5Q;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_A4 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_A5 = CLBLL_L_X42Y95_SLICE_X69Y95_BQ;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_A6 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_A4 = CLBLM_R_X41Y107_SLICE_X66Y107_DO6;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_A5 = CLBLM_R_X41Y103_SLICE_X67Y103_BO6;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_AX = CLBLL_L_X42Y95_SLICE_X69Y95_CO6;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_A6 = CLBLM_R_X41Y103_SLICE_X67Y103_CO5;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_B1 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_B2 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_B3 = CLBLL_L_X42Y93_SLICE_X68Y93_C_XOR;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_B4 = CLBLL_L_X42Y95_SLICE_X69Y95_BQ;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_B5 = CLBLL_L_X42Y96_SLICE_X68Y96_AO5;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_B6 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_B1 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_B2 = CLBLL_L_X42Y106_SLICE_X68Y106_CO5;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_C1 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_C2 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_C3 = CLBLL_L_X42Y96_SLICE_X68Y96_AO5;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_C4 = CLBLL_L_X42Y95_SLICE_X69Y95_A5Q;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_C5 = CLBLL_L_X42Y95_SLICE_X68Y95_A_XOR;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_C6 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_C1 = CLBLM_R_X41Y106_SLICE_X66Y106_BO6;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_C2 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_C3 = CLBLM_R_X41Y105_SLICE_X67Y105_AO6;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_C4 = CLBLM_R_X41Y105_SLICE_X66Y105_CO6;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_C5 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_CE = CLBLL_L_X42Y110_SLICE_X68Y110_BO6;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_D1 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_D2 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_D3 = CLBLL_L_X42Y96_SLICE_X68Y96_AO5;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_D4 = CLBLL_L_X42Y95_SLICE_X69Y95_DQ;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_D5 = CLBLL_L_X42Y94_SLICE_X68Y94_D_XOR;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_D6 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_D1 = CLBLL_L_X42Y109_SLICE_X69Y109_BO5;
  assign CLBLL_L_X42Y95_SLICE_X69Y95_DX = CLBLL_L_X42Y95_SLICE_X69Y95_DQ;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_D2 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_D3 = CLBLM_R_X41Y103_SLICE_X67Y103_D5Q;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_D4 = CLBLM_R_X41Y116_SLICE_X67Y116_DO5;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_A1 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_A2 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_A3 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_A4 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_A5 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_A6 = 1'b1;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_D1 = CLBLM_R_X3Y59_SLICE_X3Y59_B5Q;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_B1 = CLBLL_L_X42Y110_SLICE_X68Y110_AO5;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_B2 = CLBLM_R_X41Y114_SLICE_X67Y114_A5Q;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_B3 = CLBLM_R_X41Y111_SLICE_X66Y111_DQ;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_B4 = CLBLM_R_X41Y109_SLICE_X67Y109_CO5;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_A1 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_A2 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_A3 = CLBLL_L_X42Y69_SLICE_X68Y69_AO5;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_A4 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_A5 = CLBLL_L_X42Y69_SLICE_X68Y69_AQ;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_A6 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_B5 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_B6 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_AX = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_B1 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_B2 = CLBLL_L_X42Y69_SLICE_X68Y69_CQ;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_B3 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_B4 = CLBLL_L_X42Y70_SLICE_X68Y70_B_XOR;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_B5 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_B6 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_C1 = CLBLL_L_X42Y109_SLICE_X69Y109_BO5;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_C2 = CLBLM_R_X41Y109_SLICE_X67Y109_BO5;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_BX = 1'b0;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_C4 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_C1 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_C2 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_C3 = CLBLL_L_X42Y69_SLICE_X68Y69_B_XOR;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_C4 = CLBLL_L_X42Y71_SLICE_X68Y71_B5Q;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_C5 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_C6 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_D1 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_D2 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_D3 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_D4 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_D5 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_CX = 1'b0;
  assign CLBLM_R_X41Y103_SLICE_X66Y103_D6 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_D1 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_D2 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_D3 = CLBLL_L_X42Y70_SLICE_X68Y70_A_XOR;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_D4 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_D5 = CLBLL_L_X42Y70_SLICE_X68Y70_DQ;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_D6 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_DX = 1'b0;
  assign CLBLL_L_X42Y69_SLICE_X68Y69_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_A1 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_A2 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_A3 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_A4 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_A5 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_A6 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_B1 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_B2 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_B3 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_B4 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_B5 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_B6 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_C1 = CLBLL_L_X42Y69_SLICE_X68Y69_BQ;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_C2 = CLBLL_L_X42Y71_SLICE_X68Y71_B5Q;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_C3 = CLBLL_L_X42Y69_SLICE_X68Y69_DQ;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_C4 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_C5 = CLBLL_L_X42Y70_SLICE_X68Y70_DQ;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_C6 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_D1 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_D2 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_D3 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_D4 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_D5 = 1'b1;
  assign CLBLL_L_X42Y69_SLICE_X69Y69_D6 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_A1 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_A2 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_A3 = CLBLL_L_X42Y110_SLICE_X69Y110_CO6;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_A4 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_A5 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_A6 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_AX = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_B1 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_B2 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_B3 = CLBLL_L_X42Y96_SLICE_X69Y96_B5Q;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_B4 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_B5 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_B6 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_BX = 1'b0;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_C1 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_C2 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_C3 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_C4 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_C5 = CLBLL_L_X42Y96_SLICE_X69Y96_BQ;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_C6 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_CX = 1'b0;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_D1 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_D2 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_D3 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_D4 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_D5 = 1'b0;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_D6 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X68Y43_DX = 1'b0;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_A1 = CLBLL_L_X42Y96_SLICE_X68Y96_AO5;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_A2 = 1'b1;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_A3 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_A4 = CLBLL_L_X42Y92_SLICE_X68Y92_C_XOR;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_A5 = CLBLL_L_X42Y96_SLICE_X68Y96_DO6;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_A6 = 1'b1;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_AX = CLBLL_L_X42Y96_SLICE_X68Y96_BQ;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_B1 = CLBLL_L_X42Y97_SLICE_X68Y97_DO5;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_B2 = CLBLL_L_X42Y113_SLICE_X68Y113_D5Q;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_B3 = CLBLL_L_X42Y96_SLICE_X68Y96_BQ;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_B4 = 1'b1;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_B5 = CLBLL_L_X42Y93_SLICE_X68Y93_A5Q;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_B6 = 1'b1;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_BX = CLBLL_L_X42Y96_SLICE_X68Y96_CO6;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_C1 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_C2 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_C3 = CLBLL_L_X42Y96_SLICE_X68Y96_AO5;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_C4 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_A1 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_A2 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_A3 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_A4 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_A5 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_A6 = 1'b1;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_C5 = CLBLL_L_X42Y96_SLICE_X68Y96_BQ;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_C6 = 1'b1;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_B1 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_B2 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_B3 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_B4 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_B5 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_B6 = 1'b1;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_CX = CLBLL_L_X42Y96_SLICE_X68Y96_DO5;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_D1 = CLBLL_L_X42Y96_SLICE_X68Y96_CQ;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_D2 = CLBLL_L_X42Y95_SLICE_X68Y95_B_XOR;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_C1 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_C2 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_C3 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_C4 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_C5 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_C6 = 1'b1;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_DX = CLBLL_L_X42Y96_SLICE_X68Y96_CQ;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_D1 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_D2 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_D3 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_D4 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_D5 = 1'b1;
  assign CLBLL_L_X42Y43_SLICE_X69Y43_D6 = 1'b1;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_A1 = CLBLL_L_X42Y96_SLICE_X69Y96_BQ;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_A2 = CLBLL_L_X42Y112_SLICE_X69Y112_C5Q;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_A3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_A4 = CLBLL_L_X42Y71_SLICE_X68Y71_BQ;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_A5 = CLBLL_L_X42Y112_SLICE_X69Y112_DQ;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_A6 = CLBLL_L_X42Y43_SLICE_X68Y43_C_XOR;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_A1 = CLBLM_R_X41Y107_SLICE_X67Y107_BO6;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_A2 = CLBLM_R_X41Y104_SLICE_X67Y104_DO5;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_A3 = CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_B1 = 1'b1;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_B2 = CLBLL_L_X42Y96_SLICE_X69Y96_AO6;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_B3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_B4 = 1'b1;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_B5 = 1'b1;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_B6 = 1'b1;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_A4 = CLBLM_R_X41Y104_SLICE_X67Y104_DO6;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_A5 = CLBLM_R_X41Y103_SLICE_X66Y103_CO5;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_BX = CLBLL_L_X42Y71_SLICE_X68Y71_AO6;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_C1 = CLBLL_L_X42Y118_SLICE_X69Y118_B5Q;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_C2 = CLBLL_L_X42Y118_SLICE_X69Y118_A5Q;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_C3 = CLBLL_L_X42Y118_SLICE_X69Y118_CQ;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_C4 = CLBLL_L_X42Y118_SLICE_X69Y118_D5Q;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_C5 = CLBLL_L_X42Y96_SLICE_X69Y96_BQ;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_C6 = CLBLL_L_X42Y96_SLICE_X69Y96_B5Q;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_B4 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_B5 = CLBLM_R_X41Y104_SLICE_X67Y104_CO6;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_C1 = 1'b1;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_C2 = CLBLM_R_X41Y105_SLICE_X67Y105_CO6;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_C3 = CLBLM_R_X41Y105_SLICE_X67Y105_AO6;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_C4 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_D1 = CLBLL_L_X42Y96_SLICE_X69Y96_BQ;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_D2 = CLBLL_L_X42Y118_SLICE_X69Y118_DQ;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_D3 = CLBLL_L_X42Y96_SLICE_X69Y96_B5Q;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_D4 = CLBLL_L_X42Y118_SLICE_X69Y118_C5Q;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_D5 = CLBLL_L_X42Y118_SLICE_X69Y118_BQ;
  assign CLBLL_L_X42Y96_SLICE_X69Y96_D6 = CLBLL_L_X42Y118_SLICE_X69Y118_AQ;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_CX = CLBLM_R_X41Y104_SLICE_X67Y104_AO6;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_D1 = CLBLL_L_X42Y105_SLICE_X68Y105_CO5;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_D2 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_D3 = 1'b1;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_D4 = CLBLL_L_X42Y105_SLICE_X68Y105_DO6;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_D5 = 1'b1;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_D6 = 1'b1;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_A1 = CLBLM_R_X41Y107_SLICE_X67Y107_BO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_A2 = CLBLM_R_X41Y104_SLICE_X66Y104_CO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_A3 = CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_A4 = CLBLL_L_X42Y104_SLICE_X68Y104_CO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_A5 = CLBLM_R_X41Y104_SLICE_X66Y104_BO5;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_A6 = CLBLM_R_X41Y104_SLICE_X66Y104_CO5;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_A1 = CLBLL_L_X42Y69_SLICE_X68Y69_DQ;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_A2 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_A3 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_A4 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_A5 = CLBLL_L_X42Y71_SLICE_X68Y71_DO6;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_A6 = 1'b1;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_B1 = CLBLL_L_X42Y107_SLICE_X68Y107_CO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_B2 = CLBLM_R_X41Y105_SLICE_X67Y105_CO5;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_AX = 1'b0;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_B3 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_B1 = 1'b0;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_B2 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_B3 = CLBLL_L_X42Y69_SLICE_X68Y69_BQ;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_B4 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_B5 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_B6 = 1'b1;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_C3 = CLBLM_R_X41Y105_SLICE_X66Y105_AO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_C4 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_BX = CLBLL_L_X42Y71_SLICE_X68Y71_DO5;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_C5 = CLBLM_R_X41Y109_SLICE_X67Y109_AO6;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_C1 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_C2 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_C3 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_C4 = CLBLL_L_X42Y70_SLICE_X68Y70_AQ;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_C5 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_C6 = 1'b1;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_C6 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_CIN = CLBLL_L_X42Y69_SLICE_X68Y69_COUT;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_D1 = CLBLL_L_X42Y102_SLICE_X69Y102_BO5;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_D2 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_CX = 1'b0;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_D3 = CLBLM_R_X41Y100_SLICE_X67Y100_DQ;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_D1 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_D2 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_D3 = CLBLL_L_X42Y70_SLICE_X68Y70_BQ;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_D4 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_D5 = CLBLL_L_X42Y71_SLICE_X68Y71_BO6;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_D6 = 1'b1;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_D5 = 1'b1;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_D6 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X68Y70_DX = 1'b0;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_DX = CLBLM_R_X41Y104_SLICE_X66Y104_AO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_A1 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_A2 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_A3 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_A4 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_A5 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_A6 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_B1 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_B2 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_B3 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_B4 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_B5 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_B6 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_C1 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_C2 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_C3 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_C4 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_C5 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_C6 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_D1 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_D2 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_D3 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_D4 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_D5 = 1'b1;
  assign CLBLL_L_X42Y70_SLICE_X69Y70_D6 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_B5 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_D3 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_D4 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_D5 = 1'b1;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_A1 = CLBLL_L_X42Y93_SLICE_X68Y93_B_XOR;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_A2 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_A3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_A4 = CLBLL_L_X42Y96_SLICE_X68Y96_AO5;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_A5 = CLBLL_L_X42Y97_SLICE_X68Y97_BQ;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_A6 = 1'b1;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_B1 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_B2 = CLBLL_L_X42Y104_SLICE_X69Y104_BQ;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_B3 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_B4 = CLBLL_L_X42Y104_SLICE_X69Y104_AQ;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_B5 = 1'b1;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_B6 = 1'b1;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_BX = CLBLL_L_X42Y97_SLICE_X68Y97_AO5;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_C1 = CLBLL_L_X42Y113_SLICE_X68Y113_D5Q;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_C2 = CLBLL_L_X42Y92_SLICE_X69Y92_B5Q;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_C3 = CLBLL_L_X42Y97_SLICE_X68Y97_DO5;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_C4 = CLBLL_L_X42Y95_SLICE_X68Y95_D5Q;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_C5 = CLBLL_L_X42Y93_SLICE_X68Y93_A5Q;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_C6 = 1'b1;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_D1 = CLBLL_L_X42Y97_SLICE_X68Y97_BO5;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_D2 = CLBLL_L_X42Y93_SLICE_X68Y93_BQ;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_D3 = CLBLL_L_X42Y93_SLICE_X68Y93_DQ;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_D4 = CLBLL_L_X42Y104_SLICE_X69Y104_CQ;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_D5 = CLBLL_L_X42Y93_SLICE_X68Y93_CQ;
  assign CLBLL_L_X42Y97_SLICE_X68Y97_D6 = 1'b1;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_A1 = BRAM_L_X44Y95_RAMB18_X2Y38_DO4;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_A2 = BRAM_L_X44Y95_RAMB18_X2Y38_DO10;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_A3 = BRAM_L_X44Y95_RAMB18_X2Y38_DO9;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_A4 = BRAM_L_X44Y95_RAMB18_X2Y38_DOP0;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_A5 = CLBLL_L_X42Y95_SLICE_X69Y95_CQ;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_A6 = CLBLL_L_X42Y92_SLICE_X69Y92_AQ;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_A1 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_B1 = CLBLL_L_X42Y97_SLICE_X69Y97_DO6;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_B2 = BRAM_L_X44Y95_RAMB18_X2Y38_DO5;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_B3 = 1'b1;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_B4 = CLBLL_L_X42Y93_SLICE_X69Y93_CO5;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_B5 = CLBLL_L_X42Y91_SLICE_X69Y91_D5Q;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_B6 = 1'b1;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_A2 = CLBLM_R_X41Y105_SLICE_X67Y105_DO5;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_A3 = CLBLL_L_X42Y107_SLICE_X69Y107_DQ;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_A4 = CLBLM_R_X41Y107_SLICE_X66Y107_AO6;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_C1 = CLBLL_L_X42Y97_SLICE_X69Y97_BO5;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_C2 = CLBLL_L_X42Y92_SLICE_X69Y92_B5Q;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_C3 = CLBLL_L_X42Y95_SLICE_X68Y95_D5Q;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_C4 = CLBLL_L_X42Y97_SLICE_X68Y97_BO6;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_C5 = CLBLL_L_X42Y96_SLICE_X68Y96_BO6;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_C6 = 1'b1;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_CE = CLBLL_L_X42Y97_SLICE_X68Y97_CO5;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_B4 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_B5 = CLBLL_L_X42Y108_SLICE_X69Y108_D5Q;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_B6 = 1'b1;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_C1 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_C2 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_D1 = BRAM_L_X44Y95_RAMB18_X2Y38_DO7;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_D2 = CLBLL_L_X42Y95_SLICE_X69Y95_D5Q;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_D3 = BRAM_L_X44Y95_RAMB18_X2Y38_DO2;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_D4 = CLBLL_L_X42Y95_SLICE_X69Y95_AQ;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_D5 = CLBLL_L_X42Y97_SLICE_X69Y97_AO6;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_D6 = 1'b1;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_C4 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_C5 = CLBLM_R_X41Y105_SLICE_X67Y105_AO6;
  assign CLBLL_L_X42Y97_SLICE_X69Y97_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_D1 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_D2 = CLBLM_R_X41Y109_SLICE_X66Y109_BO6;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_D3 = CLBLM_R_X41Y100_SLICE_X67Y100_A5Q;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_D4 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_D5 = CLBLL_L_X42Y109_SLICE_X69Y109_DQ;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_D6 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_B3 = CLBLM_R_X41Y116_SLICE_X66Y116_CQ;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_B4 = 1'b1;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_A1 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_A2 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_A3 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_A4 = CLBLM_R_X41Y106_SLICE_X66Y106_CO6;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_A5 = CLBLM_R_X41Y105_SLICE_X66Y105_CO6;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_A1 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_A2 = CLBLL_L_X42Y71_SLICE_X68Y71_BQ;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_A3 = CLBLL_L_X42Y112_SLICE_X69Y112_DQ;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_A4 = CLBLL_L_X42Y96_SLICE_X69Y96_B5Q;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_A5 = CLBLL_L_X42Y112_SLICE_X69Y112_C5Q;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_A6 = CLBLL_L_X42Y43_SLICE_X68Y43_B_XOR;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_A6 = CLBLM_R_X41Y106_SLICE_X66Y106_AO6;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_B1 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_B1 = CLBLL_L_X42Y71_SLICE_X68Y71_CO5;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_B2 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_B3 = CLBLL_L_X42Y69_SLICE_X68Y69_D_XOR;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_B4 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_B5 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_B6 = 1'b1;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_B2 = CLBLM_R_X41Y105_SLICE_X67Y105_AO6;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_B3 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_BX = CLBLL_L_X42Y69_SLICE_X68Y69_C_XOR;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_B5 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_D3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_C1 = CLBLL_L_X42Y70_SLICE_X68Y70_AQ;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_C2 = CLBLL_L_X42Y69_SLICE_X68Y69_C_XOR;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_C3 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_C4 = CLBLL_L_X42Y69_SLICE_X69Y69_CO5;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_C5 = CLBLL_L_X42Y70_SLICE_X68Y70_BQ;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_C6 = 1'b1;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_D4 = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_C4 = CLBLL_L_X42Y108_SLICE_X69Y108_BO5;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_D5 = CLBLL_L_X42Y96_SLICE_X68Y96_AO5;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_C6 = CLBLL_L_X42Y107_SLICE_X68Y107_BO5;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_CE = CLBLL_L_X42Y110_SLICE_X68Y110_BO6;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_D1 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_D2 = CLBLL_L_X42Y71_SLICE_X68Y71_CO5;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_D3 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_D4 = CLBLL_L_X42Y70_SLICE_X68Y70_C_XOR;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_D5 = CLBLL_L_X42Y70_SLICE_X68Y70_D_XOR;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_D6 = 1'b1;
  assign CLBLL_L_X42Y96_SLICE_X68Y96_D6 = 1'b1;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_D1 = CLBLL_L_X42Y106_SLICE_X69Y106_BO5;
  assign CLBLL_L_X42Y71_SLICE_X68Y71_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_D4 = CLBLM_R_X41Y101_SLICE_X67Y101_BO5;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_D5 = CLBLM_R_X41Y105_SLICE_X66Y105_BO6;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_D6 = CLBLM_R_X41Y100_SLICE_X67Y100_BO5;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_C4 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_C5 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_A1 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_A2 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_A3 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_A4 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_A5 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_A6 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_B1 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_B2 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_B3 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_B4 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_B5 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_B6 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_C1 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_C2 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_C3 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_C4 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_C5 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_C6 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_D1 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_D2 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_D3 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_D4 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_D5 = 1'b1;
  assign CLBLL_L_X42Y71_SLICE_X69Y71_D6 = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_D1 = CLBLM_R_X3Y60_SLICE_X3Y60_B5Q;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_D5 = CLBLM_R_X41Y116_SLICE_X66Y116_D5Q;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_D6 = 1'b1;
  assign LIOI3_X0Y59_OLOGIC_X0Y59_T1 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_DX = 1'b0;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_A1 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_A2 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_A3 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_A4 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_A5 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_A6 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_B1 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_B2 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_B3 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_B4 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_B5 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_B6 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_C1 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_C2 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_C3 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_C4 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_C5 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_C6 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_D1 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_D2 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_D3 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_D4 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_D5 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X68Y98_D6 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_A1 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_A2 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_A3 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_A4 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_A5 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_A6 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_B1 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_B2 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_B3 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_B4 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_B5 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_B6 = 1'b1;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_A1 = 1'b1;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_A2 = CLBLM_R_X41Y94_SLICE_X67Y94_CQ;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_BX = BRAM_L_X44Y95_RAMB18_X2Y38_DO8;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_A3 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_C1 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_C2 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_C3 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_C4 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_C5 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_C6 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_CE = CLBLL_L_X42Y97_SLICE_X69Y97_CO6;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_A5 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_AX = CLBLM_R_X41Y114_SLICE_X66Y114_D5Q;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_B1 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_B2 = 1'b1;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_B3 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_B4 = CLBLM_R_X41Y106_SLICE_X67Y106_DO5;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_D1 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_D2 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_D3 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_D4 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_D5 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_D6 = 1'b1;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_BX = CLBLM_R_X41Y93_SLICE_X67Y93_DQ;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_C1 = 1'b1;
  assign CLBLL_L_X42Y98_SLICE_X69Y98_DX = BRAM_L_X44Y95_RAMB18_X2Y38_DO6;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_C2 = 1'b1;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_C3 = 1'b1;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_C4 = CLBLM_R_X41Y94_SLICE_X67Y94_BQ;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_C5 = 1'b1;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_C6 = 1'b1;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_CE = CLBLM_R_X41Y116_SLICE_X66Y116_DO6;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_CX = CLBLM_R_X41Y94_SLICE_X67Y94_DQ;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_D1 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_D2 = CLBLM_R_X41Y108_SLICE_X67Y108_CO6;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_D3 = CLBLM_R_X41Y106_SLICE_X67Y106_CQ;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_D4 = CLBLL_L_X42Y111_SLICE_X69Y111_DQ;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_D5 = CLBLL_L_X42Y106_SLICE_X69Y106_CO6;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_D6 = 1'b1;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_A1 = CLBLM_R_X41Y106_SLICE_X67Y106_BQ;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_A2 = CLBLL_L_X42Y107_SLICE_X68Y107_BO5;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_A3 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_A4 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_A5 = CLBLM_R_X41Y106_SLICE_X66Y106_DO5;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_A6 = CLBLM_R_X41Y107_SLICE_X66Y107_CO6;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_B1 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_B2 = CLBLM_R_X41Y106_SLICE_X66Y106_DO5;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_B3 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_B4 = CLBLM_R_X41Y106_SLICE_X67Y106_BQ;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_B5 = CLBLL_L_X42Y107_SLICE_X68Y107_BO5;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_B6 = CLBLM_R_X41Y106_SLICE_X66Y106_CO6;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_C1 = CLBLM_R_X41Y107_SLICE_X66Y107_AO6;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_C2 = CLBLM_R_X41Y100_SLICE_X67Y100_CQ;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_C3 = CLBLM_R_X41Y108_SLICE_X66Y108_CO6;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_C4 = CLBLL_L_X42Y107_SLICE_X69Y107_D5Q;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_C5 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_C6 = CLBLL_L_X42Y106_SLICE_X68Y106_BO5;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_D1 = CLBLL_L_X42Y107_SLICE_X69Y107_BQ;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_D2 = CLBLL_L_X42Y108_SLICE_X68Y108_BO5;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_D3 = CLBLM_R_X41Y107_SLICE_X66Y107_AO6;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_D4 = CLBLM_R_X41Y108_SLICE_X66Y108_CO6;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_D5 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLM_R_X41Y106_SLICE_X66Y106_D6 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_D5 = CLBLL_L_X42Y97_SLICE_X69Y97_C5Q;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_D6 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_DX = CLBLM_R_X41Y114_SLICE_X66Y114_BO6;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_A6 = CLBLM_R_X41Y104_SLICE_X67Y104_BO5;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_B1 = CLBLL_L_X42Y105_SLICE_X68Y105_CO6;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_B2 = CLBLL_L_X42Y103_SLICE_X68Y103_AO6;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_B3 = CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_B6 = 1'b1;
  assign CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_CE0 = 1'b1;
  assign CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_CE1 = 1'b1;
  assign CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_IGNORE0 = 1'b1;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_A1 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_A2 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_A3 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_A4 = CLBLM_R_X41Y107_SLICE_X66Y107_BO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_A5 = CLBLM_R_X41Y107_SLICE_X67Y107_BO5;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_A6 = CLBLM_R_X41Y106_SLICE_X66Y106_BO6;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_C5 = CLBLL_L_X42Y107_SLICE_X68Y107_AO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_B1 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_C6 = 1'b1;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_B2 = CLBLL_L_X42Y103_SLICE_X69Y103_BQ;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_B3 = 1'b1;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_B4 = CLBLM_R_X41Y107_SLICE_X66Y107_CO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_B5 = CLBLL_L_X42Y109_SLICE_X69Y109_CO5;
  assign CLBLM_R_X41Y104_SLICE_X67Y104_CE = CLBLL_L_X42Y110_SLICE_X68Y110_BO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_B6 = 1'b1;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_C1 = CLBLM_R_X41Y107_SLICE_X67Y107_DO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_C2 = CLBLM_R_X41Y111_SLICE_X66Y111_BO5;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_C3 = CLBLM_R_X41Y107_SLICE_X67Y107_AO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_C4 = CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_C5 = CLBLM_R_X41Y107_SLICE_X67Y107_BO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_C6 = CLBLM_R_X41Y101_SLICE_X66Y101_BO5;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_CE = CLBLL_L_X42Y110_SLICE_X68Y110_BO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_D1 = 1'b1;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_D2 = CLBLL_L_X42Y111_SLICE_X69Y111_CO5;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_D3 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_D4 = CLBLM_R_X41Y110_SLICE_X67Y110_CO5;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_D5 = CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_D6 = 1'b1;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_DX = CLBLM_R_X41Y107_SLICE_X67Y107_CO6;
  assign CLBLM_R_X41Y107_SLICE_X67Y107_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_A1 = CLBLM_R_X41Y108_SLICE_X66Y108_D5Q;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_A2 = CLBLM_R_X41Y109_SLICE_X66Y109_AQ;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_A3 = CLBLL_L_X42Y109_SLICE_X68Y109_DQ;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_A4 = CLBLM_R_X41Y108_SLICE_X67Y108_CO5;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_A5 = CLBLL_L_X42Y106_SLICE_X69Y106_CO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_A6 = CLBLM_R_X41Y108_SLICE_X67Y108_DO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_B1 = CLBLL_L_X42Y68_SLICE_X68Y68_BQ;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_B2 = CLBLL_L_X42Y108_SLICE_X68Y108_AO5;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_B3 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_B4 = CLBLM_R_X41Y107_SLICE_X66Y107_AO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_B5 = CLBLM_R_X41Y108_SLICE_X66Y108_CO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_B6 = CLBLL_L_X42Y107_SLICE_X68Y107_BO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_C1 = CLBLM_R_X41Y108_SLICE_X66Y108_CO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_C2 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_C3 = CLBLM_R_X41Y107_SLICE_X66Y107_AO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_C4 = CLBLL_L_X42Y107_SLICE_X69Y107_B5Q;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_C5 = CLBLM_R_X41Y106_SLICE_X67Y106_A5Q;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_C6 = CLBLL_L_X42Y108_SLICE_X68Y108_DO5;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_D1 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_D2 = CLBLM_R_X41Y106_SLICE_X67Y106_BO5;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_D3 = CLBLM_R_X41Y107_SLICE_X66Y107_BO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_D4 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_D5 = CLBLM_R_X41Y101_SLICE_X67Y101_DO6;
  assign CLBLM_R_X41Y107_SLICE_X66Y107_D6 = CLBLM_R_X41Y107_SLICE_X67Y107_BO5;
  assign LIOB33_X0Y55_IOB_X0Y55_O = CLBLM_R_X3Y59_SLICE_X3Y59_B5Q;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_B4 = CLBLM_R_X41Y105_SLICE_X67Y105_CO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_B5 = CLBLM_R_X41Y104_SLICE_X66Y104_DO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_B6 = 1'b1;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_C1 = CLBLM_R_X41Y109_SLICE_X67Y109_DO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_C2 = CLBLL_L_X42Y109_SLICE_X69Y109_BO5;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_CE = CLBLM_R_X41Y101_SLICE_X66Y101_DO5;
  assign CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_I0 = RIOB33_X57Y125_IOB_X1Y126_I;
  assign CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_I1 = 1'b1;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_A1 = CLBLM_R_X41Y115_SLICE_X66Y115_DO6;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_A2 = CLBLL_L_X42Y110_SLICE_X69Y110_BO6;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_A3 = CLBLL_L_X42Y109_SLICE_X68Y109_DO6;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_A4 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_A5 = CLBLM_R_X41Y108_SLICE_X67Y108_D5Q;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_A6 = CLBLM_R_X41Y110_SLICE_X66Y110_DO5;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_B1 = CLBLM_R_X41Y109_SLICE_X66Y109_AQ;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_B2 = CLBLM_R_X41Y108_SLICE_X67Y108_CO5;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_B3 = CLBLM_R_X41Y108_SLICE_X66Y108_D5Q;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_B4 = CLBLL_L_X42Y109_SLICE_X68Y109_DQ;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_B5 = CLBLM_R_X41Y108_SLICE_X67Y108_CO6;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_B6 = CLBLM_R_X41Y108_SLICE_X67Y108_DO6;
  assign CLBLM_R_X41Y104_SLICE_X66Y104_D4 = CLBLL_L_X42Y107_SLICE_X68Y107_BO5;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_C1 = CLBLM_R_X41Y109_SLICE_X67Y109_D5Q;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_C2 = CLBLM_R_X41Y108_SLICE_X67Y108_D5Q;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_C3 = CLBLL_L_X42Y108_SLICE_X68Y108_C5Q;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_C4 = CLBLM_R_X41Y102_SLICE_X67Y102_C5Q;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_C5 = CLBLL_L_X42Y109_SLICE_X69Y109_DQ;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_C6 = 1'b1;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_D1 = 1'b1;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_D2 = CLBLM_R_X41Y110_SLICE_X66Y110_B5Q;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_D3 = CLBLL_L_X42Y109_SLICE_X68Y109_D5Q;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_D4 = CLBLL_L_X42Y102_SLICE_X68Y102_BQ;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_D5 = 1'b1;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_D6 = 1'b1;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_DX = CLBLM_R_X41Y108_SLICE_X67Y108_AO6;
  assign CLBLM_R_X41Y108_SLICE_X67Y108_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_A1 = CLBLL_L_X42Y109_SLICE_X68Y109_DO6;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_A2 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_A3 = CLBLM_R_X41Y115_SLICE_X66Y115_DO6;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_A4 = CLBLL_L_X42Y109_SLICE_X68Y109_DQ;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_A5 = CLBLM_R_X41Y108_SLICE_X66Y108_CO5;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_A6 = CLBLM_R_X41Y110_SLICE_X66Y110_CO6;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_B1 = CLBLM_R_X41Y111_SLICE_X66Y111_AQ;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_B2 = CLBLM_R_X41Y108_SLICE_X66Y108_CO5;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_B3 = CLBLM_R_X41Y107_SLICE_X67Y107_D5Q;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_B4 = CLBLM_R_X41Y114_SLICE_X67Y114_B5Q;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_B5 = CLBLL_L_X42Y110_SLICE_X69Y110_BO5;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_B6 = CLBLM_R_X41Y110_SLICE_X66Y110_DO5;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_C1 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_C2 = CLBLM_R_X41Y108_SLICE_X67Y108_CO5;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_C3 = CLBLL_L_X42Y109_SLICE_X68Y109_DQ;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_C4 = CLBLL_L_X42Y109_SLICE_X68Y109_BO6;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_C5 = CLBLM_R_X41Y108_SLICE_X66Y108_D5Q;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_C6 = 1'b1;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_CE = CLBLM_R_X41Y108_SLICE_X66Y108_DO6;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_D1 = CLBLM_R_X41Y108_SLICE_X66Y108_CO5;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_D2 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_D3 = CLBLM_R_X41Y115_SLICE_X66Y115_DO6;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_D4 = CLBLL_L_X42Y109_SLICE_X68Y109_DO6;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_D5 = 1'b1;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_D6 = 1'b1;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_DX = CLBLM_R_X41Y108_SLICE_X66Y108_CO5;
  assign CLBLM_R_X41Y108_SLICE_X66Y108_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign LIOB33_X0Y57_IOB_X0Y57_O = CLBLM_R_X3Y60_SLICE_X3Y60_BQ;
  assign LIOI3_X0Y55_OLOGIC_X0Y55_T1 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_A1 = CLBLL_L_X42Y96_SLICE_X69Y96_DO6;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_A2 = CLBLL_L_X42Y110_SLICE_X69Y110_C5Q;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_A3 = CLBLL_L_X42Y112_SLICE_X69Y112_C5Q;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_A4 = CLBLL_L_X42Y96_SLICE_X69Y96_CO6;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_A5 = CLBLL_L_X42Y112_SLICE_X69Y112_DQ;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_A6 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_B1 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_B2 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_B3 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_B4 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_B5 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_B6 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_C1 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_C2 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_C3 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_C4 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_C5 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_C6 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_CE = CLBLL_L_X42Y71_SLICE_X68Y71_BQ;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_D1 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_D2 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_D3 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_D4 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_D5 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_D6 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X68Y101_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_A1 = BRAM_L_X44Y95_RAMB18_X2Y38_DO11;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_A2 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_A3 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_A4 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_A5 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_A6 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_AX = CLBLL_L_X42Y95_SLICE_X69Y95_D5Q;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_B1 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_B2 = CLBLM_R_X41Y111_SLICE_X66Y111_BQ;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_B3 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_B4 = CLBLL_L_X42Y106_SLICE_X69Y106_CO5;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_B5 = CLBLL_L_X42Y68_SLICE_X68Y68_C5Q;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_B6 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_BX = CLBLL_L_X42Y95_SLICE_X69Y95_CQ;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_C1 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_C2 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_C3 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_C4 = CLBLL_L_X42Y91_SLICE_X69Y91_AQ;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_C5 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_C6 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_CE = CLBLL_L_X42Y97_SLICE_X69Y97_CO6;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_A1 = CLBLL_L_X42Y68_SLICE_X68Y68_AQ;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_A2 = CLBLL_L_X42Y110_SLICE_X68Y110_AO5;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_A3 = CLBLM_R_X41Y114_SLICE_X67Y114_CQ;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_A4 = CLBLM_R_X41Y109_SLICE_X67Y109_BO6;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_CX = CLBLL_L_X42Y91_SLICE_X69Y91_D5Q;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_A5 = CLBLM_R_X41Y109_SLICE_X67Y109_CO5;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_D1 = CLBLL_L_X42Y107_SLICE_X68Y107_BO5;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_D2 = CLBLL_L_X42Y106_SLICE_X69Y106_CO5;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_D3 = CLBLL_L_X42Y68_SLICE_X68Y68_A5Q;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_D4 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_D5 = CLBLM_R_X41Y95_SLICE_X67Y95_BQ;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_D6 = 1'b1;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_A6 = 1'b1;
  assign CLBLL_L_X42Y101_SLICE_X69Y101_DX = CLBLL_L_X42Y95_SLICE_X69Y95_AQ;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_B1 = CLBLM_R_X41Y108_SLICE_X66Y108_D5Q;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_B2 = CLBLM_R_X41Y109_SLICE_X67Y109_D5Q;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_B3 = CLBLL_L_X42Y109_SLICE_X68Y109_DQ;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_B4 = CLBLM_R_X41Y108_SLICE_X67Y108_D5Q;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_B5 = CLBLL_L_X42Y109_SLICE_X68Y109_BO6;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_B6 = 1'b1;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_C1 = CLBLL_L_X42Y109_SLICE_X68Y109_DQ;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_C2 = CLBLM_R_X41Y108_SLICE_X67Y108_CO5;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_C3 = 1'b1;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_C4 = CLBLM_R_X41Y108_SLICE_X66Y108_D5Q;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_C5 = CLBLL_L_X42Y109_SLICE_X68Y109_BO6;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_C6 = 1'b1;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_CE = CLBLL_L_X42Y109_SLICE_X68Y109_DO6;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_IGNORE1 = 1'b1;
  assign CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_S0 = 1'b1;
  assign CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_S1 = 1'b1;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_D1 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_D2 = CLBLM_R_X41Y110_SLICE_X66Y110_CO6;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_D3 = CLBLM_R_X41Y102_SLICE_X66Y102_BQ;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_D4 = CLBLM_R_X41Y104_SLICE_X66Y104_D5Q;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_D5 = CLBLM_R_X41Y109_SLICE_X66Y109_CO5;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_D6 = 1'b1;
  assign CLBLM_R_X41Y109_SLICE_X67Y109_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_A1 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_A2 = CLBLM_R_X41Y102_SLICE_X66Y102_BQ;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_A3 = CLBLM_R_X41Y109_SLICE_X66Y109_CO6;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_A4 = CLBLM_R_X41Y109_SLICE_X66Y109_CO5;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_A5 = CLBLM_R_X41Y115_SLICE_X66Y115_BQ;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_A6 = 1'b1;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_B1 = CLBLM_R_X41Y109_SLICE_X67Y109_CO6;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_B2 = CLBLL_L_X42Y108_SLICE_X68Y108_C5Q;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_B3 = CLBLM_R_X41Y102_SLICE_X67Y102_C5Q;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_B4 = 1'b1;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_B5 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_B6 = 1'b1;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_C1 = CLBLL_L_X42Y102_SLICE_X68Y102_BQ;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_C2 = CLBLM_R_X41Y110_SLICE_X66Y110_B5Q;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_C3 = CLBLM_R_X41Y109_SLICE_X66Y109_AQ;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_C4 = CLBLL_L_X42Y109_SLICE_X68Y109_D5Q;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_C5 = CLBLM_R_X41Y109_SLICE_X66Y109_DO5;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_C6 = 1'b1;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_CE = CLBLL_L_X42Y109_SLICE_X68Y109_DO6;
  assign LIOB33_X0Y59_IOB_X0Y59_O = CLBLM_R_X3Y60_SLICE_X3Y60_B5Q;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_D1 = CLBLL_L_X42Y109_SLICE_X68Y109_DQ;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_D2 = CLBLM_R_X41Y108_SLICE_X66Y108_D5Q;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_D3 = CLBLM_R_X41Y108_SLICE_X67Y108_CO5;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_D4 = CLBLL_L_X42Y109_SLICE_X69Y109_DQ;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_D5 = CLBLM_R_X41Y109_SLICE_X66Y109_BO6;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_D6 = 1'b1;
  assign CLBLM_R_X41Y109_SLICE_X66Y109_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_D5 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_A1 = CLBLL_L_X42Y102_SLICE_X68Y102_DO6;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_A2 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_A3 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_A4 = CLBLL_L_X42Y103_SLICE_X69Y103_B_XOR;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_A5 = CLBLL_L_X42Y103_SLICE_X69Y103_AO5;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_A6 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_B1 = CLBLL_L_X42Y102_SLICE_X68Y102_AO6;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_B2 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_B3 = CLBLM_R_X41Y102_SLICE_X66Y102_CO6;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_B4 = CLBLL_L_X42Y110_SLICE_X69Y110_BO6;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_B5 = CLBLM_R_X41Y107_SLICE_X67Y107_D5Q;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_B6 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_C1 = CLBLM_R_X41Y102_SLICE_X66Y102_BO5;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_C2 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_C3 = CLBLM_R_X41Y102_SLICE_X66Y102_CO6;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_C4 = CLBLM_R_X41Y109_SLICE_X67Y109_CO6;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_C5 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_C6 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_CE = CLBLL_L_X42Y102_SLICE_X68Y102_DO5;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_D1 = CLBLL_L_X42Y102_SLICE_X68Y102_CO5;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_D2 = CLBLL_L_X42Y109_SLICE_X69Y109_CO6;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_D3 = CLBLL_L_X42Y103_SLICE_X68Y103_CO6;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_D4 = CLBLM_R_X41Y115_SLICE_X66Y115_DO6;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_D5 = CLBLM_R_X41Y107_SLICE_X66Y107_AO6;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_D6 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X68Y102_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_A1 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_A2 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_A3 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_A4 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_A5 = CLBLL_L_X42Y112_SLICE_X68Y112_DQ;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_A6 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_AX = CLBLL_L_X42Y112_SLICE_X68Y112_D5Q;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_B1 = CLBLL_L_X42Y106_SLICE_X69Y106_CO5;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_B2 = CLBLL_L_X42Y102_SLICE_X69Y102_D5Q;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_B3 = CLBLL_L_X42Y102_SLICE_X69Y102_DQ;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_B4 = CLBLL_L_X42Y102_SLICE_X69Y102_A5Q;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_B5 = CLBLL_L_X42Y102_SLICE_X68Y102_CO6;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_B6 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_C1 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_C2 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_C3 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_C4 = CLBLL_L_X42Y112_SLICE_X68Y112_BQ;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_C5 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_C6 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_CE = CLBLM_R_X41Y114_SLICE_X66Y114_DO6;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_CX = CLBLL_L_X42Y113_SLICE_X69Y113_A5Q;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_A1 = CLBLM_R_X41Y107_SLICE_X67Y107_BO6;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_D1 = CLBLL_L_X42Y111_SLICE_X68Y111_B5Q;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_D2 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_D3 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_D4 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_D5 = 1'b1;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_D6 = 1'b1;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_A2 = CLBLM_R_X41Y110_SLICE_X67Y110_CO5;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_A3 = CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  assign CLBLL_L_X42Y102_SLICE_X69Y102_DX = CLBLL_L_X42Y101_SLICE_X69Y101_D5Q;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_A4 = CLBLL_L_X42Y111_SLICE_X69Y111_CO5;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_A5 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_A6 = CLBLM_R_X41Y110_SLICE_X67Y110_DO5;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_B1 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_B2 = CLBLL_L_X42Y110_SLICE_X68Y110_DO6;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_B3 = CLBLM_R_X41Y110_SLICE_X67Y110_B5Q;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_B4 = CLBLM_R_X41Y110_SLICE_X67Y110_AO6;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_B5 = CLBLM_R_X41Y111_SLICE_X66Y111_CO5;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_B6 = 1'b1;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_C1 = CLBLL_L_X42Y101_SLICE_X69Y101_DO6;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_C2 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_C3 = CLBLL_L_X42Y106_SLICE_X68Y106_CO5;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_C4 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_C5 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_C6 = 1'b1;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_CE = CLBLL_L_X42Y110_SLICE_X68Y110_BO6;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_D1 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_D2 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_D3 = CLBLM_R_X41Y107_SLICE_X66Y107_BO6;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_D4 = CLBLM_R_X41Y107_SLICE_X67Y107_BO5;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_D5 = CLBLM_R_X41Y106_SLICE_X66Y106_BO6;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_D6 = 1'b1;
  assign CLBLM_R_X41Y110_SLICE_X67Y110_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_A1 = CLBLM_R_X41Y115_SLICE_X66Y115_DO6;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_A2 = CLBLM_R_X41Y110_SLICE_X66Y110_B5Q;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_A3 = CLBLM_R_X41Y110_SLICE_X66Y110_DO5;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_A4 = CLBLM_R_X41Y109_SLICE_X66Y109_AQ;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_A5 = CLBLL_L_X42Y109_SLICE_X68Y109_DO6;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_A6 = 1'b1;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_B1 = CLBLM_R_X41Y110_SLICE_X66Y110_DO6;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_B2 = CLBLM_R_X41Y109_SLICE_X66Y109_CO5;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_B3 = CLBLL_L_X42Y109_SLICE_X69Y109_BO5;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_B4 = 1'b1;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_B5 = CLBLM_R_X41Y109_SLICE_X66Y109_CO6;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_B6 = 1'b1;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_C1 = CLBLM_R_X41Y109_SLICE_X67Y109_D5Q;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_C2 = CLBLL_L_X42Y109_SLICE_X68Y109_DQ;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_C3 = CLBLL_L_X42Y109_SLICE_X68Y109_BO6;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_C4 = CLBLM_R_X41Y108_SLICE_X66Y108_D5Q;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_C5 = CLBLM_R_X41Y108_SLICE_X67Y108_D5Q;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_C6 = 1'b1;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_CE = CLBLM_R_X41Y110_SLICE_X66Y110_AO5;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_D1 = CLBLM_R_X41Y110_SLICE_X66Y110_CO5;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_D2 = 1'b1;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_D3 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_D4 = CLBLL_L_X42Y110_SLICE_X69Y110_BO6;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_D5 = CLBLM_R_X41Y110_SLICE_X66Y110_CO6;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_D6 = 1'b1;
  assign CLBLM_R_X41Y110_SLICE_X66Y110_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_A1 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_A2 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_A3 = CLBLM_R_X3Y54_SLICE_X3Y54_B5Q;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_A4 = CLBLM_R_X3Y54_SLICE_X3Y54_AO5;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_A5 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_A6 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_AX = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_B1 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_B2 = CLBLM_R_X3Y54_SLICE_X3Y54_AO5;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_B3 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_B4 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_B5 = CLBLM_R_X3Y54_SLICE_X3Y54_BQ;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_B6 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_BX = 1'b0;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_C1 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_C2 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_C3 = CLBLM_R_X3Y54_SLICE_X3Y54_CQ;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_C4 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_C5 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_C6 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_CX = 1'b0;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_D1 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_D2 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_D3 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_D4 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_D5 = CLBLM_R_X3Y54_SLICE_X3Y54_DQ;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_D6 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X3Y54_DX = 1'b0;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_A1 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_A2 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_A3 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_A4 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_A5 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_A6 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_B1 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_B2 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_B3 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_B4 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_B5 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_B6 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_C1 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_C2 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_C3 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_C4 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_C5 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_C6 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_D1 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_D2 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_D3 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_D4 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_D5 = 1'b1;
  assign CLBLM_R_X3Y54_SLICE_X2Y54_D6 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_A1 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_A2 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_A3 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_A4 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_A5 = CLBLM_R_X41Y106_SLICE_X66Y106_CO6;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_A6 = CLBLM_R_X41Y105_SLICE_X66Y105_CO6;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_B1 = CLBLL_L_X42Y103_SLICE_X68Y103_CQ;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_B2 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_B3 = CLBLL_L_X42Y103_SLICE_X68Y103_DQ;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_B4 = CLBLL_L_X42Y103_SLICE_X68Y103_BQ;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_B5 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_B6 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_BX = CLBLL_L_X42Y104_SLICE_X69Y104_BO5;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_C1 = CLBLL_L_X42Y102_SLICE_X68Y102_DO6;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_C2 = CLBLL_L_X42Y102_SLICE_X68Y102_AO6;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_C3 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_C4 = CLBLM_R_X41Y108_SLICE_X67Y108_BO6;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_C5 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_C6 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_CE = CLBLL_L_X42Y103_SLICE_X68Y103_DO5;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_CX = CLBLL_L_X42Y104_SLICE_X69Y104_CO5;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_D1 = CLBLL_L_X42Y109_SLICE_X69Y109_BO5;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_D2 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_D3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_D4 = CLBLL_L_X42Y103_SLICE_X68Y103_CO5;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_D5 = CLBLM_R_X41Y109_SLICE_X66Y109_BO5;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_D6 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X68Y103_DX = CLBLL_L_X42Y104_SLICE_X69Y104_DO5;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_A1 = CLBLL_L_X42Y103_SLICE_X69Y103_C_XOR;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_A2 = CLBLL_L_X42Y104_SLICE_X69Y104_A_XOR;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_A3 = CLBLL_L_X42Y104_SLICE_X68Y104_DO5;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_A4 = CLBLL_L_X42Y103_SLICE_X69Y103_D_XOR;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_A5 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_A6 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_AX = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_B1 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_B2 = CLBLL_L_X42Y103_SLICE_X69Y103_B_XOR;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_B3 = CLBLL_L_X42Y103_SLICE_X69Y103_BQ;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_B4 = CLBLL_L_X42Y110_SLICE_X68Y110_BO5;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_B5 = CLBLM_R_X41Y108_SLICE_X67Y108_BO6;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_B6 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_BX = 1'b0;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_C1 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_C2 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_C3 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_C4 = CLBLL_L_X42Y103_SLICE_X68Y103_DQ;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_C5 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_C6 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_CE = CLBLL_L_X42Y103_SLICE_X68Y103_DO5;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_CX = 1'b0;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_D1 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_D2 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_D3 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_D4 = 1'b1;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_D5 = CLBLL_L_X42Y103_SLICE_X68Y103_CQ;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_D6 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_A1 = CLBLL_L_X42Y109_SLICE_X69Y109_BO5;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_A2 = CLBLL_L_X42Y105_SLICE_X68Y105_AO6;
  assign CLBLL_L_X42Y103_SLICE_X69Y103_DX = 1'b0;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_A3 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_A4 = CLBLM_R_X41Y111_SLICE_X67Y111_A5Q;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_A5 = CLBLM_R_X41Y111_SLICE_X67Y111_BO5;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_A6 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_B1 = CLBLM_R_X41Y108_SLICE_X66Y108_CO5;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_B2 = CLBLM_R_X41Y115_SLICE_X67Y115_BQ;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_B3 = CLBLL_L_X42Y110_SLICE_X69Y110_BO5;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_B4 = CLBLL_L_X42Y102_SLICE_X69Y102_CQ;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_B5 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_B6 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_C1 = CLBLM_R_X41Y108_SLICE_X66Y108_CO5;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_C2 = CLBLM_R_X41Y106_SLICE_X67Y106_AQ;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_C3 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_C4 = CLBLL_L_X42Y102_SLICE_X69Y102_AQ;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_C5 = CLBLL_L_X42Y110_SLICE_X69Y110_BO5;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_C6 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_CE = CLBLL_L_X42Y110_SLICE_X68Y110_BO6;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_D1 = CLBLM_R_X41Y105_SLICE_X66Y105_DQ;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_D2 = CLBLL_L_X42Y109_SLICE_X69Y109_BO5;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_D3 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_D4 = CLBLM_R_X41Y110_SLICE_X66Y110_DO6;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_D5 = CLBLM_R_X41Y111_SLICE_X67Y111_CO5;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_D6 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X67Y111_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_A1 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_A2 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_A3 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_A4 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_A5 = CLBLL_L_X42Y113_SLICE_X69Y113_BQ;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_A6 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_AX = CLBLL_L_X42Y113_SLICE_X69Y113_D5Q;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_B1 = CLBLM_R_X41Y109_SLICE_X67Y109_BO6;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_B2 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_B3 = CLBLL_L_X42Y102_SLICE_X68Y102_BO5;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_B4 = CLBLL_L_X42Y109_SLICE_X69Y109_BO5;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_B5 = CLBLM_R_X41Y108_SLICE_X66Y108_BO6;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_B6 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_BX = CLBLL_L_X42Y113_SLICE_X69Y113_B5Q;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_C1 = CLBLL_L_X42Y110_SLICE_X68Y110_AO5;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_C2 = CLBLM_R_X41Y115_SLICE_X67Y115_AQ;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_C3 = CLBLM_R_X41Y111_SLICE_X66Y111_A5Q;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_C4 = CLBLM_R_X41Y111_SLICE_X66Y111_DO5;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_C5 = CLBLM_R_X41Y109_SLICE_X67Y109_CO5;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_C6 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_CE = CLBLM_R_X41Y114_SLICE_X66Y114_DO6;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_D1 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_D2 = CLBLL_L_X42Y110_SLICE_X68Y110_DO6;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_D3 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_D4 = CLBLL_L_X42Y109_SLICE_X69Y109_BO5;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_D5 = CLBLM_R_X41Y110_SLICE_X67Y110_B5Q;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_D6 = 1'b1;
  assign CLBLM_R_X41Y111_SLICE_X66Y111_DX = CLBLL_L_X42Y113_SLICE_X69Y113_DQ;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_A1 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_A2 = CLBLM_R_X3Y55_SLICE_X3Y55_B5Q;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_A3 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_A4 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_A5 = CLBLM_R_X3Y55_SLICE_X3Y55_D_XOR;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_A6 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_AX = 1'b0;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_B1 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_B2 = CLBLM_R_X3Y55_SLICE_X3Y55_BQ;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_B3 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_B4 = CLBLM_R_X3Y55_SLICE_X3Y55_A_XOR;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_B5 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_B6 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_BX = 1'b0;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_C1 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_C2 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_C3 = CLBLM_R_X3Y55_SLICE_X3Y55_DQ;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_C4 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_C5 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_C6 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_CIN = CLBLM_R_X3Y54_SLICE_X3Y54_COUT;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_A6 = CLBLM_R_X41Y105_SLICE_X67Y105_BO5;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_CX = 1'b0;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_D1 = CLBLM_R_X3Y55_SLICE_X3Y55_C_XOR;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_D2 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_D3 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_D4 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_D5 = CLBLM_R_X3Y55_SLICE_X3Y55_AQ;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_D6 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X3Y55_DX = 1'b0;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_A1 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_A2 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_A3 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_A4 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_A5 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_A6 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_B1 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_B2 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_B3 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_B4 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_B5 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_B6 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_C1 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_C2 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_C3 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_C4 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_C5 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_C6 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_D1 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_D2 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_D3 = 1'b1;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_A1 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_A2 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_A3 = CLBLL_L_X42Y106_SLICE_X68Y106_DO5;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_A4 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_A5 = CLBLL_L_X42Y105_SLICE_X68Y105_BO5;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_A6 = CLBLL_L_X42Y101_SLICE_X69Y101_DO6;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_D4 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_D5 = 1'b1;
  assign CLBLM_R_X3Y55_SLICE_X2Y55_D6 = 1'b1;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_B1 = CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_B2 = CLBLL_L_X42Y104_SLICE_X68Y104_AO6;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_B3 = CLBLM_R_X41Y107_SLICE_X67Y107_BO6;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_B4 = CLBLL_L_X42Y104_SLICE_X68Y104_DO6;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_B5 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_B6 = CLBLM_R_X41Y105_SLICE_X66Y105_AO6;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_C1 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_C2 = CLBLM_R_X41Y106_SLICE_X67Y106_BO6;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_C3 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_C4 = CLBLL_L_X42Y105_SLICE_X69Y105_BO6;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_C5 = CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_C6 = CLBLL_L_X42Y104_SLICE_X68Y104_AO6;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_CE = CLBLL_L_X42Y103_SLICE_X68Y103_DO5;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_A5 = CLBLM_R_X41Y108_SLICE_X66Y108_CO6;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR0 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR1 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR2 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR3 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR4 = CLBLL_L_X42Y94_SLICE_X68Y94_BQ;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR5 = CLBLL_L_X42Y90_SLICE_X68Y90_BQ;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR6 = CLBLL_L_X42Y90_SLICE_X68Y90_DQ;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_D1 = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR9 = CLBLL_L_X42Y91_SLICE_X68Y91_BQ;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR10 = CLBLL_L_X42Y91_SLICE_X68Y91_CQ;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_D2 = CLBLL_L_X42Y105_SLICE_X69Y105_BO6;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_D3 = CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR13 = CLBLL_L_X42Y92_SLICE_X69Y92_DQ;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRATIEHIGH0 = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRATIEHIGH1 = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBTIEHIGH0 = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBTIEHIGH1 = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR0 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR1 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR2 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR3 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR4 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR5 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR6 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR7 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR8 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR9 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR10 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR11 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR12 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRBWRADDR13 = 1'b0;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_B1 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_B2 = CLBLL_L_X42Y107_SLICE_X69Y107_CQ;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_RDCLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_WRCLK = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI0 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI1 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI2 = 1'b0;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_A3 = CLBLL_L_X42Y103_SLICE_X68Y103_BQ;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI3 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI4 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI5 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI6 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI7 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI8 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI9 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI10 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI11 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI12 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI13 = 1'b0;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_A6 = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI0 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI1 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI2 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI3 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI4 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI5 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI6 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI7 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI8 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI9 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI10 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI11 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI12 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI13 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI14 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIBDI15 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIPADIP0 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIPADIP1 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIPBDIP0 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIPBDIP1 = 1'b0;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_D1 = CLBLL_L_X42Y103_SLICE_X68Y103_DQ;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_D2 = CLBLL_L_X42Y110_SLICE_X68Y110_BO5;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_D3 = CLBLM_R_X41Y108_SLICE_X67Y108_BO6;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_D4 = 1'b0;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_D5 = CLBLL_L_X42Y103_SLICE_X69Y103_C_XOR;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_D6 = 1'b1;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_CX = 1'b0;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_DX = 1'b0;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_B3 = CLBLM_R_X41Y108_SLICE_X67Y108_BO6;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_C3 = CLBLL_L_X42Y107_SLICE_X68Y107_AO6;
  assign CLBLM_R_X41Y105_SLICE_X67Y105_C6 = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_RDEN = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_WREN = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_REGCE = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_REGCEB = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_RDRCLK = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_REGCLKB = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_RST = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_RSTRAMB = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_RSTREG = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_RSTREGB = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_WEA0 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_WEA1 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_WEA2 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_WEA3 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE0 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE1 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE2 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE3 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE4 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE5 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE6 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_WEBWE7 = 1'b0;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_A1 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_A2 = CLBLM_R_X3Y56_SLICE_X3Y56_B5Q;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_A3 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_A4 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_A5 = CLBLM_R_X3Y56_SLICE_X3Y56_D_XOR;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_A6 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_AX = 1'b0;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_B1 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_B2 = CLBLM_R_X3Y56_SLICE_X3Y56_BQ;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_B3 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_B4 = CLBLM_R_X3Y56_SLICE_X3Y56_A_XOR;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_B5 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_B6 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_BX = 1'b0;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_C1 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_C2 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_C3 = CLBLM_R_X3Y56_SLICE_X3Y56_DQ;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_C4 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_C5 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_C6 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_CIN = CLBLM_R_X3Y55_SLICE_X3Y55_COUT;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_CX = 1'b0;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_D1 = CLBLM_R_X3Y56_SLICE_X3Y56_C_XOR;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_D2 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_D3 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_D4 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_D5 = CLBLM_R_X3Y56_SLICE_X3Y56_AQ;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_D6 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X3Y56_DX = 1'b0;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_A1 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_A2 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_A3 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_A4 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_A5 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_A6 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_B1 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_B2 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_B3 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_B4 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_B5 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_B6 = 1'b1;
  assign LIOI3_X0Y67_OLOGIC_X0Y68_D1 = CLBLM_R_X3Y59_SLICE_X3Y59_AQ;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_C1 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_C2 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_C3 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_C4 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_C5 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_C6 = 1'b1;
  assign LIOI3_X0Y67_OLOGIC_X0Y68_T1 = 1'b1;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_A1 = CLBLM_R_X41Y101_SLICE_X67Y101_C5Q;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_A2 = CLBLL_L_X42Y105_SLICE_X68Y105_CO5;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_A3 = CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_A4 = CLBLM_R_X41Y107_SLICE_X67Y107_BO6;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_A5 = CLBLL_L_X42Y105_SLICE_X68Y105_DO6;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_A6 = CLBLL_L_X42Y105_SLICE_X68Y105_CO6;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_D1 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_D2 = 1'b1;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_B1 = CLBLL_L_X42Y105_SLICE_X68Y105_CQ;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_B2 = CLBLM_R_X41Y114_SLICE_X67Y114_DQ;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_B3 = CLBLL_L_X42Y106_SLICE_X69Y106_DO5;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_B4 = CLBLL_L_X42Y107_SLICE_X68Y107_BO5;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_B5 = CLBLL_L_X42Y106_SLICE_X69Y106_CO5;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_B6 = 1'b1;
  assign CLBLM_R_X3Y56_SLICE_X2Y56_D6 = 1'b1;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_B4 = CLBLM_R_X41Y105_SLICE_X66Y105_CO6;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_C1 = CLBLL_L_X42Y105_SLICE_X68Y105_BO5;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_C2 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_C3 = CLBLM_R_X41Y106_SLICE_X67Y106_BO6;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_C4 = 1'b1;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_C5 = CLBLM_R_X41Y106_SLICE_X66Y106_AO6;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_C6 = 1'b1;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_CE = CLBLM_R_X41Y114_SLICE_X66Y114_DO6;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_B6 = CLBLM_R_X41Y106_SLICE_X66Y106_BO6;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_CX = CLBLL_L_X42Y92_SLICE_X68Y92_CQ;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_D1 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_D2 = CLBLL_L_X42Y106_SLICE_X68Y106_DO5;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_D3 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_D4 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_D5 = CLBLL_L_X42Y105_SLICE_X69Y105_BO6;
  assign CLBLL_L_X42Y105_SLICE_X68Y105_D6 = CLBLL_L_X42Y101_SLICE_X69Y101_DO6;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_D1 = CLBLM_R_X3Y60_SLICE_X3Y60_BQ;
  assign LIOI3_TBYTESRC_X0Y57_OLOGIC_X0Y57_T1 = 1'b1;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_C1 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_C2 = CLBLM_R_X41Y100_SLICE_X67Y100_C5Q;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_C3 = CLBLM_R_X41Y108_SLICE_X66Y108_CO6;
  assign LIOB33_X0Y67_IOB_X0Y68_O = CLBLM_R_X3Y59_SLICE_X3Y59_AQ;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_A1 = 1'b1;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_A2 = 1'b1;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_A3 = CLBLL_L_X42Y101_SLICE_X69Y101_A5Q;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_A4 = 1'b1;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_A5 = 1'b1;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_A6 = 1'b1;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_C5 = CLBLL_L_X42Y102_SLICE_X69Y102_C5Q;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_AX = CLBLL_L_X42Y101_SLICE_X69Y101_AQ;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_C3 = CLBLM_R_X41Y93_SLICE_X67Y93_BQ;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_B1 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_B2 = CLBLL_L_X42Y106_SLICE_X68Y106_DO5;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_B3 = CLBLL_L_X42Y105_SLICE_X69Y105_CO5;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_B4 = CLBLL_L_X42Y105_SLICE_X69Y105_DO5;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_B5 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_B6 = 1'b1;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_C1 = CLBLL_L_X42Y105_SLICE_X69Y105_A5Q;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_C2 = CLBLM_R_X41Y95_SLICE_X67Y95_CQ;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_C3 = CLBLL_L_X42Y106_SLICE_X69Y106_CO6;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_C4 = CLBLM_R_X41Y108_SLICE_X67Y108_CO6;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_C5 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_C6 = 1'b1;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_CE = CLBLM_R_X41Y114_SLICE_X66Y114_DO6;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_C6 = 1'b1;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_I = CLK_BUFG_TOP_R_X78Y105_BUFGCTRL_X0Y16_O;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_D1 = CLBLM_R_X41Y108_SLICE_X67Y108_CO6;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_D2 = CLBLM_R_X41Y95_SLICE_X67Y95_DQ;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_D3 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_D4 = CLBLL_L_X42Y106_SLICE_X69Y106_CO6;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_D5 = CLBLL_L_X42Y111_SLICE_X69Y111_D5Q;
  assign CLBLL_L_X42Y105_SLICE_X69Y105_D6 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_D2 = CLBLM_R_X41Y111_SLICE_X67Y111_DO5;
  assign CLBLM_R_X41Y105_SLICE_X66Y105_D3 = CLBLM_R_X41Y107_SLICE_X67Y107_BO6;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_D5 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_D6 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X67Y100_DX = CLBLM_R_X41Y92_SLICE_X67Y92_CQ;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_A3 = 1'b1;
  assign CLBLM_R_X41Y100_SLICE_X66Y100_A4 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_AX = 1'b0;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_A1 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_A2 = CLBLM_R_X3Y57_SLICE_X3Y57_DQ;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_A3 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_A4 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_A5 = CLBLM_R_X3Y57_SLICE_X3Y57_C_XOR;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_A6 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_AX = 1'b0;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_B1 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_B2 = CLBLM_R_X3Y57_SLICE_X3Y57_BQ;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_B3 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_B4 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_B5 = CLBLM_R_X3Y57_SLICE_X3Y57_D_XOR;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_B6 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_BX = 1'b0;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_C1 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_C2 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_C3 = CLBLM_R_X3Y57_SLICE_X3Y57_AQ;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_C4 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_C5 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_C6 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_CIN = CLBLM_R_X3Y56_SLICE_X3Y56_COUT;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_CX = 1'b0;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_D1 = CLBLM_R_X3Y57_SLICE_X3Y57_A_XOR;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_D2 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_D3 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_D4 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_D5 = CLBLM_R_X3Y57_SLICE_X3Y57_B5Q;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_D6 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X3Y57_DX = 1'b0;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_A1 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_A2 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_A3 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_A4 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_A5 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_A6 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_B1 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_B2 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_B3 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_B4 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_B5 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_B6 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_C1 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_C2 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_C3 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_C4 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_C5 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_C6 = 1'b1;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_A1 = 1'b1;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_A2 = 1'b1;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_A3 = 1'b1;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_A4 = 1'b1;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_A5 = CLBLL_L_X42Y98_SLICE_X69Y98_D5Q;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_A6 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_D1 = 1'b1;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_AX = CLBLL_L_X42Y113_SLICE_X69Y113_CQ;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_D2 = 1'b1;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_B1 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_B2 = CLBLL_L_X42Y109_SLICE_X69Y109_BO6;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_D6 = 1'b1;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_B3 = CLBLL_L_X42Y106_SLICE_X68Y106_AQ;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_B4 = CLBLL_L_X42Y106_SLICE_X68Y106_A5Q;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_B5 = CLBLL_L_X42Y108_SLICE_X68Y108_C5Q;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_B6 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_D3 = 1'b1;
  assign CLBLM_R_X3Y57_SLICE_X2Y57_D4 = 1'b1;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_C1 = CLBLL_L_X42Y106_SLICE_X69Y106_CO5;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_C2 = CLBLM_R_X41Y114_SLICE_X67Y114_DQ;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_C3 = CLBLL_L_X42Y105_SLICE_X68Y105_CQ;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_C4 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_C5 = CLBLM_R_X41Y107_SLICE_X66Y107_AO6;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_C6 = 1'b1;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_CE = CLBLM_R_X41Y114_SLICE_X66Y114_DO6;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_D1 = CLBLL_L_X42Y106_SLICE_X69Y106_CO6;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_D2 = CLBLL_L_X42Y107_SLICE_X69Y107_C5Q;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_D3 = CLBLM_R_X41Y95_SLICE_X67Y95_AQ;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_D4 = CLBLM_R_X41Y108_SLICE_X67Y108_CO6;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_D5 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLL_L_X42Y106_SLICE_X68Y106_D6 = 1'b1;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_A1 = CLBLL_L_X42Y106_SLICE_X69Y106_DO5;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_A2 = CLBLL_L_X42Y108_SLICE_X69Y108_AQ;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_A3 = CLBLM_R_X41Y108_SLICE_X66Y108_CO6;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_A4 = CLBLM_R_X41Y100_SLICE_X67Y100_AQ;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_A5 = CLBLL_L_X42Y107_SLICE_X68Y107_BO5;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_A6 = CLBLL_L_X42Y106_SLICE_X69Y106_DO6;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_B1 = CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_B2 = CLBLM_R_X41Y105_SLICE_X67Y105_CO6;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_B3 = CLBLL_L_X42Y106_SLICE_X69Y106_AO6;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_B4 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_B5 = CLBLL_L_X42Y107_SLICE_X68Y107_CO6;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_B6 = 1'b1;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_C1 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_C2 = CLBLM_R_X41Y102_SLICE_X67Y102_C5Q;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_C3 = 1'b1;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_C4 = CLBLL_L_X42Y109_SLICE_X69Y109_DQ;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_C5 = CLBLL_L_X42Y108_SLICE_X68Y108_C5Q;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_C6 = 1'b1;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_CE = CLBLM_R_X41Y114_SLICE_X66Y114_DO6;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_CX = CLBLL_L_X42Y80_SLICE_X69Y80_B5Q;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_D1 = CLBLL_L_X42Y106_SLICE_X69Y106_CQ;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_D2 = CLBLL_L_X42Y68_SLICE_X68Y68_CQ;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_D3 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_D4 = CLBLL_L_X42Y106_SLICE_X69Y106_CO5;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_D5 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLL_L_X42Y106_SLICE_X69Y106_D6 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_A1 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_A2 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_A3 = CLBLM_R_X41Y114_SLICE_X66Y114_BO5;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_A4 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_A5 = CLBLM_R_X41Y116_SLICE_X66Y116_D5Q;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_A6 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_A1 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_A2 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_A3 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_A4 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_A5 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_A6 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_AX = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_B1 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_B2 = CLBLM_R_X41Y114_SLICE_X66Y114_DQ;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_B1 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_B2 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_B3 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_B4 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_B5 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_B6 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_B6 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_BX = 1'b0;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_C1 = CLBLM_R_X41Y114_SLICE_X66Y114_DQ;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_C1 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_C2 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_C3 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_C4 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_C5 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_C6 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_C6 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_CE = CLBLM_R_X41Y116_SLICE_X66Y116_DO6;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_CX = 1'b0;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_D1 = CLBLM_R_X41Y93_SLICE_X67Y93_C5Q;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_D2 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_D3 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X67Y114_D4 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_D1 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_D2 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_D3 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_D4 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_D5 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X68Y80_D6 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_A1 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_A2 = CLBLM_R_X41Y114_SLICE_X66Y114_DQ;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_A3 = CLBLM_R_X41Y115_SLICE_X66Y115_BO5;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_A4 = CLBLL_L_X42Y97_SLICE_X69Y97_C5Q;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_A5 = CLBLM_R_X41Y114_SLICE_X66Y114_D5Q;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_A6 = CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_B1 = CLBLM_R_X41Y115_SLICE_X66Y115_BO5;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_B2 = CLBLM_R_X41Y114_SLICE_X66Y114_D5Q;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_B3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_B4 = CLBLL_L_X42Y97_SLICE_X69Y97_C5Q;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_B5 = CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_B6 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_C1 = CLBLL_L_X42Y97_SLICE_X69Y97_C5Q;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_C2 = CLBLM_R_X41Y115_SLICE_X67Y115_D_XOR;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_C3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_C4 = CLBLM_R_X41Y114_SLICE_X66Y114_CQ;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_C5 = CLBLM_R_X41Y115_SLICE_X66Y115_BO5;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_C6 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_A1 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_A2 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_A3 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_A4 = BRAM_L_X44Y95_RAMB18_X2Y38_DO3;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_A5 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_A6 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_AX = CLBLL_L_X42Y96_SLICE_X68Y96_DQ;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_D1 = CLBLM_R_X41Y114_SLICE_X66Y114_AO6;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_B1 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_B2 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_B3 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_B4 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_B5 = BRAM_L_X44Y95_RAMB18_X2Y38_DO1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_B6 = 1'b1;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_D2 = CLBLM_R_X41Y102_SLICE_X66Y102_BQ;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_D3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_BX = BRAM_L_X44Y95_RAMB18_X2Y38_DO0;
  assign CLBLM_R_X41Y114_SLICE_X66Y114_D4 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_C1 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_C2 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_C3 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_C4 = BRAM_L_X44Y95_RAMB18_X2Y38_DO13;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_C5 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_C6 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_CE = CLBLL_L_X42Y97_SLICE_X69Y97_CO6;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_CX = CLBLL_L_X42Y92_SLICE_X69Y92_DQ;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_A1 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_D1 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_D2 = CLBLL_L_X42Y96_SLICE_X68Y96_AQ;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_A4 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_A5 = CLBLM_R_X3Y58_SLICE_X3Y58_C_XOR;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_A6 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_D3 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_D4 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_D5 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_D6 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_A2 = CLBLM_R_X3Y58_SLICE_X3Y58_DQ;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_A3 = 1'b1;
  assign CLBLL_L_X42Y80_SLICE_X69Y80_DX = CLBLL_L_X42Y93_SLICE_X68Y93_A5Q;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_B1 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_B2 = CLBLM_R_X3Y58_SLICE_X3Y58_BQ;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_B3 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_B4 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_B5 = CLBLM_R_X3Y58_SLICE_X3Y58_D_XOR;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_B6 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_BX = 1'b0;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_C1 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_C2 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_C3 = CLBLM_R_X3Y58_SLICE_X3Y58_AQ;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_C4 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_C5 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_C6 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_CIN = CLBLM_R_X3Y57_SLICE_X3Y57_COUT;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_CX = 1'b0;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_D1 = CLBLM_R_X3Y58_SLICE_X3Y58_A_XOR;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_D2 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_D3 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_D4 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_D5 = CLBLM_R_X3Y58_SLICE_X3Y58_B5Q;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_D6 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X3Y58_DX = 1'b0;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_A1 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_A2 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_A3 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_A4 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_A5 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_A6 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_B1 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_B2 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_B3 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_B4 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_B5 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_B6 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_C1 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_C2 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_C3 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_C4 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_A1 = CLBLM_R_X41Y108_SLICE_X66Y108_CO6;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_A2 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_A3 = CLBLL_L_X42Y107_SLICE_X68Y107_DO5;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_A4 = CLBLM_R_X41Y100_SLICE_X67Y100_BQ;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_A5 = CLBLL_L_X42Y107_SLICE_X69Y107_A5Q;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_A6 = CLBLL_L_X42Y107_SLICE_X68Y107_BO5;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_C5 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_C6 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_B1 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_B2 = CLBLM_R_X41Y107_SLICE_X66Y107_AO6;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_B3 = CLBLM_R_X41Y106_SLICE_X67Y106_C5Q;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_B4 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_D3 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_B5 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_B6 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_D1 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_BX = CLBLL_L_X42Y101_SLICE_X69Y101_C5Q;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_D2 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_C1 = CLBLM_R_X41Y100_SLICE_X67Y100_D5Q;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_C2 = CLBLL_L_X42Y107_SLICE_X68Y107_BO5;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_C3 = CLBLL_L_X42Y103_SLICE_X68Y103_BO5;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_C4 = CLBLM_R_X41Y108_SLICE_X66Y108_CO6;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_C5 = CLBLL_L_X42Y107_SLICE_X69Y107_AQ;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_C6 = CLBLL_L_X42Y101_SLICE_X69Y101_BO5;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_CE = CLBLM_R_X41Y114_SLICE_X66Y114_DO6;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_D5 = 1'b1;
  assign CLBLM_R_X3Y58_SLICE_X2Y58_D6 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_D1 = CLBLL_L_X42Y68_SLICE_X68Y68_DQ;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_D2 = CLBLM_R_X41Y108_SLICE_X67Y108_BO6;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_D3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_D4 = CLBLL_L_X42Y107_SLICE_X68Y107_BQ;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_D5 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLL_L_X42Y107_SLICE_X68Y107_D6 = 1'b1;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_C6 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_A1 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_A2 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_A3 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_A4 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_A5 = CLBLL_L_X42Y112_SLICE_X68Y112_B5Q;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_A6 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_AX = CLBLL_L_X42Y112_SLICE_X68Y112_C5Q;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_B1 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_B2 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_B3 = CLBLL_L_X42Y92_SLICE_X68Y92_D5Q;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_B4 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_B5 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_B6 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_BX = CLBLL_L_X42Y112_SLICE_X68Y112_CQ;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_C1 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_C2 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_C3 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_C4 = CLBLL_L_X42Y92_SLICE_X68Y92_AQ;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_C5 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_C6 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_CE = CLBLM_R_X41Y114_SLICE_X66Y114_DO6;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_CX = CLBLL_L_X42Y92_SLICE_X68Y92_BQ;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_D1 = CLBLL_L_X42Y112_SLICE_X68Y112_AQ;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_D2 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_D3 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_D4 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_D5 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_D6 = 1'b1;
  assign CLBLL_L_X42Y107_SLICE_X69Y107_DX = CLBLL_L_X42Y112_SLICE_X68Y112_A5Q;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_A1 = CLBLM_R_X41Y115_SLICE_X66Y115_DQ;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_A2 = CLBLM_R_X41Y115_SLICE_X66Y115_D5Q;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_A3 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_A4 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_A5 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_A6 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_AX = 1'b0;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_B1 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_B2 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_B3 = CLBLM_R_X41Y114_SLICE_X66Y114_CQ;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_B4 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_B5 = CLBLM_R_X41Y116_SLICE_X66Y116_DQ;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_B6 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_BX = 1'b0;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_C1 = CLBLM_R_X41Y115_SLICE_X66Y115_DQ;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_C2 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_C3 = CLBLM_R_X41Y115_SLICE_X66Y115_D5Q;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_C4 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_C5 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_C6 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_CE = CLBLM_R_X41Y116_SLICE_X66Y116_DO6;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_CIN = CLBLM_R_X41Y114_SLICE_X67Y114_COUT;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_CX = 1'b0;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_D1 = CLBLM_R_X41Y114_SLICE_X66Y114_CQ;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_D2 = CLBLM_R_X41Y116_SLICE_X66Y116_DQ;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_D3 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_D4 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_D5 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_D6 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X67Y115_DX = 1'b0;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_A1 = CLBLM_R_X41Y115_SLICE_X66Y115_BO5;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_A2 = CLBLM_R_X41Y115_SLICE_X66Y115_DQ;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_A3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_A4 = CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_A5 = CLBLL_L_X42Y97_SLICE_X69Y97_C5Q;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_A6 = CLBLM_R_X41Y115_SLICE_X67Y115_A_XOR;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_B1 = CLBLM_R_X41Y115_SLICE_X66Y115_BQ;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_B2 = CLBLM_R_X41Y107_SLICE_X66Y107_AO6;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_B3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_B4 = CLBLL_L_X42Y103_SLICE_X68Y103_CO6;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_B5 = CLBLL_L_X42Y90_SLICE_X69Y90_CQ;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_B6 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_C1 = CLBLM_R_X41Y115_SLICE_X66Y115_BO5;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_C2 = CLBLL_L_X42Y97_SLICE_X69Y97_C5Q;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_C3 = CLBLM_R_X41Y115_SLICE_X66Y115_D5Q;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_C4 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_C5 = CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_C6 = CLBLM_R_X41Y115_SLICE_X67Y115_C_XOR;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_D1 = CLBLM_R_X41Y109_SLICE_X66Y109_CO5;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_D2 = CLBLM_R_X41Y115_SLICE_X66Y115_BQ;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_D3 = CLBLM_R_X41Y115_SLICE_X66Y115_AO6;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_D4 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_D5 = CLBLM_R_X41Y102_SLICE_X66Y102_BQ;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_D6 = 1'b1;
  assign CLBLM_R_X41Y115_SLICE_X66Y115_DX = CLBLM_R_X41Y115_SLICE_X66Y115_CO6;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_A1 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_A2 = CLBLM_R_X3Y59_SLICE_X3Y59_DQ;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_A3 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_A4 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_A5 = CLBLM_R_X3Y59_SLICE_X3Y59_C_XOR;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_A6 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_AX = 1'b0;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_B1 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_B2 = CLBLM_R_X3Y59_SLICE_X3Y59_BQ;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_B3 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_B4 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_B5 = CLBLM_R_X3Y59_SLICE_X3Y59_D_XOR;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_B6 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_BX = 1'b0;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_C1 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_C2 = CLBLM_R_X3Y59_SLICE_X3Y59_AQ;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_C3 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_C4 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_C5 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_C6 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_CIN = CLBLM_R_X3Y58_SLICE_X3Y58_COUT;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_CX = 1'b0;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_D1 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_D2 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_D3 = CLBLM_R_X3Y59_SLICE_X3Y59_B5Q;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_D4 = CLBLM_R_X3Y59_SLICE_X3Y59_A_XOR;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_D5 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_D6 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X3Y59_DX = 1'b0;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_A1 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_A2 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_A3 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_A4 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_A5 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_A6 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_B1 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_B2 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_B3 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_B4 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_B5 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_B6 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_A1 = CLBLL_L_X42Y108_SLICE_X68Y108_C5Q;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_A2 = CLBLL_L_X42Y109_SLICE_X69Y109_BO6;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_A3 = CLBLL_L_X42Y68_SLICE_X68Y68_D5Q;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_A4 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_A5 = CLBLL_L_X42Y111_SLICE_X69Y111_BQ;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_A6 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_C1 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_C2 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_C3 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_B1 = CLBLL_L_X42Y105_SLICE_X69Y105_AQ;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_B2 = CLBLL_L_X42Y111_SLICE_X69Y111_AQ;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_B3 = CLBLL_L_X42Y109_SLICE_X69Y109_BO6;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_B4 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_B5 = CLBLL_L_X42Y108_SLICE_X68Y108_C5Q;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_B6 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_D1 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_D2 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_C1 = CLBLL_L_X42Y102_SLICE_X68Y102_AO6;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_C2 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_C3 = CLBLL_L_X42Y109_SLICE_X69Y109_CO6;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_C4 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_C5 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_C6 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_CE = CLBLM_R_X41Y102_SLICE_X66Y102_AO5;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_D3 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_D4 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_D5 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_D6 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_D1 = CLBLL_L_X42Y107_SLICE_X68Y107_DO6;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_D2 = CLBLL_L_X42Y108_SLICE_X68Y108_C5Q;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_D3 = CLBLL_L_X42Y68_SLICE_X68Y68_B5Q;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_D4 = CLBLL_L_X42Y111_SLICE_X69Y111_A5Q;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_D5 = CLBLL_L_X42Y109_SLICE_X69Y109_BO6;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_D6 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X68Y108_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_A1 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_A2 = CLBLL_L_X42Y111_SLICE_X68Y111_DQ;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_A3 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_A4 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_A5 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_A6 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_AX = CLBLL_L_X42Y111_SLICE_X68Y111_D5Q;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_B1 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_B2 = CLBLL_L_X42Y108_SLICE_X69Y108_DQ;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_B3 = CLBLM_R_X41Y108_SLICE_X67Y108_BO6;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_B4 = CLBLL_L_X42Y108_SLICE_X69Y108_A5Q;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_B5 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_B6 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_C1 = CLBLM_R_X41Y102_SLICE_X66Y102_AO6;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_C2 = CLBLM_R_X41Y108_SLICE_X67Y108_BO6;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_C3 = CLBLL_L_X42Y102_SLICE_X68Y102_AO5;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_C4 = CLBLL_L_X42Y104_SLICE_X68Y104_DQ;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_C5 = CLBLL_L_X42Y110_SLICE_X68Y110_BO5;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_C6 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_CE = CLBLM_R_X41Y114_SLICE_X66Y114_DO6;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_D5 = CLBLM_R_X41Y103_SLICE_X67Y103_AO6;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_D1 = CLBLL_L_X42Y111_SLICE_X68Y111_C5Q;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_D2 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_D3 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_D4 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_D5 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_D6 = 1'b1;
  assign CLBLL_L_X42Y108_SLICE_X69Y108_DX = CLBLL_L_X42Y101_SLICE_X69Y101_CQ;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_D6 = 1'b1;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_A1 = 1'b0;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_A2 = 1'b1;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_A3 = 1'b1;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_A4 = 1'b1;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_A5 = CLBLL_L_X42Y113_SLICE_X69Y113_AQ;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_A6 = 1'b1;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_AX = 1'b0;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_B1 = CLBLM_R_X41Y109_SLICE_X67Y109_CO5;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_B2 = CLBLM_R_X41Y115_SLICE_X67Y115_DQ;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_B3 = 1'b0;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_B4 = CLBLM_R_X41Y116_SLICE_X67Y116_AQ;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_B5 = CLBLL_L_X42Y110_SLICE_X68Y110_AO5;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_B6 = 1'b1;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_BX = 1'b0;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_C1 = 1'b1;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_C2 = CLBLL_L_X42Y113_SLICE_X69Y113_C5Q;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_C3 = 1'b1;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_C4 = 1'b0;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_C5 = 1'b1;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_C6 = 1'b1;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_CE = CLBLM_R_X41Y114_SLICE_X66Y114_DO6;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_CIN = CLBLM_R_X41Y115_SLICE_X67Y115_COUT;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_CX = 1'b0;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_D1 = CLBLM_R_X41Y109_SLICE_X67Y109_CO5;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_D2 = CLBLM_R_X41Y116_SLICE_X67Y116_CQ;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_D3 = CLBLM_R_X41Y115_SLICE_X67Y115_CQ;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_D4 = 1'b0;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_D5 = CLBLL_L_X42Y110_SLICE_X68Y110_AO5;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_D6 = 1'b1;
  assign CLBLM_R_X41Y116_SLICE_X67Y116_DX = 1'b0;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_A1 = CLBLM_R_X41Y115_SLICE_X66Y115_BO5;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_A2 = CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_A3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_A4 = CLBLL_L_X42Y97_SLICE_X69Y97_C5Q;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_A5 = CLBLM_R_X41Y116_SLICE_X66Y116_DQ;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_A6 = CLBLM_R_X41Y115_SLICE_X67Y115_B_XOR;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_B1 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_B2 = CLBLM_R_X41Y116_SLICE_X66Y116_D5Q;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_B3 = CLBLM_R_X41Y115_SLICE_X66Y115_BO5;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_B4 = CLBLM_R_X41Y114_SLICE_X67Y114_D_XOR;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_B5 = CLBLL_L_X42Y97_SLICE_X69Y97_C5Q;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_B6 = CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_C1 = CLBLM_R_X41Y116_SLICE_X66Y116_CQ;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_C2 = CLBLM_R_X41Y115_SLICE_X66Y115_BO5;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_C3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_C4 = CLBLM_R_X41Y114_SLICE_X67Y114_C_XOR;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_C5 = CLBLL_L_X42Y97_SLICE_X69Y97_C5Q;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_C6 = CLBLM_R_X41Y116_SLICE_X67Y116_A_XOR;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLM_R_X41Y103_SLICE_X67Y103_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_D1 = 1'b1;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_D2 = 1'b1;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_D3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_D4 = CLBLM_R_X41Y115_SLICE_X66Y115_BO5;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_D5 = CLBLM_R_X41Y116_SLICE_X66Y116_AO6;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_D6 = 1'b1;
  assign CLBLM_R_X41Y116_SLICE_X66Y116_DX = CLBLM_R_X41Y116_SLICE_X66Y116_BO6;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_A1 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_A2 = CLBLM_R_X3Y60_SLICE_X3Y60_B5Q;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_A3 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_A4 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_A5 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_A6 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_AX = 1'b0;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_B1 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_B2 = CLBLM_R_X3Y60_SLICE_X3Y60_BQ;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_B3 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_B4 = CLBLM_R_X3Y60_SLICE_X3Y60_A_XOR;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_B5 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_B6 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_BX = 1'b0;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_C1 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_C2 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_C3 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_C4 = 1'b0;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_C5 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_C6 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_CIN = CLBLM_R_X3Y59_SLICE_X3Y59_COUT;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X0Y20_O;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_CX = 1'b0;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_D1 = 1'b0;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_D2 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_D3 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_D4 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_D5 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_D6 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X3Y60_DX = 1'b0;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_A1 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_A2 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_A3 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_A4 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_A5 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_A6 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_B1 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_B2 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_B3 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_B4 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_B5 = 1'b1;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_A1 = CLBLL_L_X42Y110_SLICE_X69Y110_BO5;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_A2 = CLBLL_L_X42Y109_SLICE_X68Y109_DO6;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_A3 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_A4 = CLBLM_R_X41Y115_SLICE_X66Y115_DO6;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_A5 = CLBLL_L_X42Y109_SLICE_X68Y109_D5Q;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_C1 = 1'b1;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_A6 = CLBLM_R_X41Y109_SLICE_X66Y109_CO6;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_C4 = 1'b1;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_B1 = CLBLM_R_X41Y102_SLICE_X67Y102_C5Q;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_C6 = 1'b1;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_B2 = CLBLL_L_X42Y108_SLICE_X68Y108_C5Q;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_B3 = CLBLL_L_X42Y109_SLICE_X69Y109_DQ;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_B4 = CLBLL_L_X42Y102_SLICE_X68Y102_BQ;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_B5 = CLBLL_L_X42Y109_SLICE_X68Y109_D5Q;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_B6 = CLBLM_R_X41Y110_SLICE_X66Y110_AO6;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_C3 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_C5 = 1'b1;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_C1 = CLBLL_L_X42Y109_SLICE_X68Y109_D5Q;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_D1 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_D2 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_D3 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_D4 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_D5 = 1'b1;
  assign CLBLM_R_X3Y60_SLICE_X2Y60_D6 = 1'b1;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_C2 = CLBLM_R_X41Y108_SLICE_X66Y108_D5Q;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_C3 = CLBLM_R_X41Y110_SLICE_X66Y110_AO6;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_C4 = CLBLL_L_X42Y102_SLICE_X68Y102_BQ;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_C5 = CLBLL_L_X42Y109_SLICE_X68Y109_DQ;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_C6 = CLBLM_R_X41Y108_SLICE_X67Y108_CO5;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_D1 = 1'b1;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_D3 = CLBLM_R_X41Y109_SLICE_X66Y109_BO5;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_D4 = 1'b1;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_D5 = CLBLM_R_X41Y102_SLICE_X66Y102_AO6;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_D6 = 1'b1;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_D2 = CLBLL_L_X42Y109_SLICE_X68Y109_AO6;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_DX = CLBLM_R_X41Y108_SLICE_X66Y108_AO6;
  assign CLBLL_L_X42Y109_SLICE_X68Y109_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_A4 = 1'b1;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_A6 = 1'b1;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_A1 = CLBLL_L_X42Y110_SLICE_X69Y110_AQ;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_A2 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_A3 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_A4 = CLBLL_L_X42Y109_SLICE_X69Y109_BO5;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_A5 = CLBLM_R_X41Y109_SLICE_X66Y109_CO6;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_A6 = CLBLL_L_X42Y110_SLICE_X68Y110_DO5;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_B1 = CLBLL_L_X42Y110_SLICE_X68Y110_AO5;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_B2 = CLBLL_L_X42Y109_SLICE_X69Y109_DQ;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_B3 = CLBLM_R_X41Y102_SLICE_X67Y102_C5Q;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_B4 = CLBLL_L_X42Y109_SLICE_X69Y109_CO5;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_B5 = CLBLM_R_X41Y109_SLICE_X67Y109_CO5;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_B6 = 1'b1;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_C1 = CLBLM_R_X41Y109_SLICE_X67Y109_CO6;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_C2 = CLBLL_L_X42Y109_SLICE_X68Y109_CO6;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_C3 = CLBLL_L_X42Y108_SLICE_X68Y108_C5Q;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_C4 = CLBLM_R_X41Y102_SLICE_X67Y102_C5Q;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_C5 = CLBLL_L_X42Y109_SLICE_X69Y109_DQ;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_C6 = 1'b1;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_CE = CLBLL_L_X42Y110_SLICE_X69Y110_AO5;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_D1 = CLBLL_L_X42Y109_SLICE_X69Y109_DQ;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_D2 = CLBLL_L_X42Y110_SLICE_X68Y110_AO5;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_D3 = CLBLM_R_X41Y102_SLICE_X66Y102_CO6;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_D4 = CLBLL_L_X42Y103_SLICE_X68Y103_CO6;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_D5 = 1'b1;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_D6 = 1'b1;
  assign CLBLL_L_X42Y109_SLICE_X69Y109_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_B5 = CLBLM_R_X41Y107_SLICE_X66Y107_BO6;
  assign CLBLM_R_X41Y106_SLICE_X67Y106_B6 = 1'b1;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_A1 = CLBLM_R_X41Y110_SLICE_X66Y110_AO6;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_A2 = CLBLL_L_X42Y102_SLICE_X68Y102_BQ;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_A3 = CLBLM_R_X41Y109_SLICE_X66Y109_DO5;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_A4 = CLBLL_L_X42Y109_SLICE_X68Y109_D5Q;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_A5 = 1'b1;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_A6 = 1'b1;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_B1 = CLBLL_L_X42Y109_SLICE_X69Y109_CO5;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_B2 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_B3 = CLBLL_L_X42Y110_SLICE_X68Y110_DO5;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_B4 = CLBLL_L_X42Y109_SLICE_X69Y109_BO5;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_B5 = CLBLM_R_X41Y109_SLICE_X66Y109_CO6;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_B6 = 1'b1;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_C1 = CLBLL_L_X42Y110_SLICE_X68Y110_C5Q;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_C2 = CLBLL_L_X42Y109_SLICE_X69Y109_BO5;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_C3 = CLBLM_R_X41Y116_SLICE_X67Y116_BO5;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_C4 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_C5 = CLBLL_L_X42Y104_SLICE_X68Y104_BO6;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_C6 = 1'b1;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_CE = CLBLL_L_X42Y110_SLICE_X68Y110_BO6;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_D1 = 1'b1;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_D2 = CLBLM_R_X41Y109_SLICE_X67Y109_BO6;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_D3 = CLBLL_L_X42Y110_SLICE_X68Y110_DO6;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_D4 = CLBLM_R_X41Y109_SLICE_X67Y109_BO5;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_D5 = CLBLL_L_X42Y110_SLICE_X68Y110_AO6;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_D6 = 1'b1;
  assign CLBLL_L_X42Y110_SLICE_X68Y110_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_A1 = CLBLL_L_X42Y109_SLICE_X68Y109_DO6;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_A2 = CLBLM_R_X41Y115_SLICE_X66Y115_DO6;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_A3 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_A4 = CLBLL_L_X42Y110_SLICE_X69Y110_BO5;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_A5 = 1'b1;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_A6 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_B5 = CLBLM_R_X41Y104_SLICE_X66Y104_DO6;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_B6 = 1'b1;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_AX = CLBLL_L_X42Y110_SLICE_X69Y110_DO5;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_B1 = CLBLM_R_X41Y109_SLICE_X66Y109_DO5;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_B2 = CLBLL_L_X42Y102_SLICE_X68Y102_BQ;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_B3 = 1'b1;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_B4 = CLBLL_L_X42Y109_SLICE_X68Y109_D5Q;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_B5 = CLBLM_R_X41Y110_SLICE_X66Y110_AO6;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_B6 = 1'b1;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_BX = CLBLL_L_X42Y109_SLICE_X69Y109_AO6;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_C1 = CLBLL_L_X42Y110_SLICE_X69Y110_C5Q;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_C2 = CLBLL_L_X42Y71_SLICE_X68Y71_BQ;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_C3 = CLBLL_L_X42Y112_SLICE_X69Y112_DQ;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_C4 = CLBLL_L_X42Y112_SLICE_X69Y112_C5Q;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_C5 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_C6 = 1'b1;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_D1 = CLBLL_L_X42Y71_SLICE_X68Y71_BQ;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_D2 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_D3 = CLBLL_L_X42Y110_SLICE_X69Y110_AQ;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_D4 = CLBLL_L_X42Y112_SLICE_X69Y112_BQ;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_D5 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLL_L_X42Y110_SLICE_X69Y110_D6 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_C3 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_C4 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_C5 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_C6 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_CE = CLBLM_R_X41Y102_SLICE_X67Y102_DO5;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_A1 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_A2 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_A3 = CLBLM_R_X41Y92_SLICE_X67Y92_BQ;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_A4 = CLBLM_R_X41Y92_SLICE_X67Y92_AO5;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_A5 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_A6 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_AX = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_B1 = CLBLM_R_X41Y92_SLICE_X67Y92_AO5;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_B2 = CLBLM_R_X41Y92_SLICE_X67Y92_DQ;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_B3 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_B4 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_B5 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_B6 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_BX = 1'b0;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_C1 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_C2 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_C3 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_C4 = CLBLM_R_X41Y92_SLICE_X67Y92_CQ;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_C5 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_C6 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_CE = CLBLL_L_X42Y90_SLICE_X69Y90_CQ;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_CX = 1'b0;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_D1 = CLBLM_R_X41Y94_SLICE_X67Y94_B5Q;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_D2 = CLBLM_R_X41Y92_SLICE_X67Y92_B_XOR;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_D3 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_D4 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_D5 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_D6 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_DX = 1'b0;
  assign CLBLM_R_X41Y92_SLICE_X67Y92_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_A1 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_A2 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_A3 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_A4 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_A5 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_A6 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_D6 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_B1 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_B2 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_B3 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_B4 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_B5 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_B6 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_C1 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_C2 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_C3 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_C4 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_C5 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_C6 = 1'b1;
  assign CLBLM_R_X41Y101_SLICE_X67Y101_DX = CLBLM_R_X41Y101_SLICE_X67Y101_CO6;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_D1 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_D2 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_D3 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_D4 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_D5 = 1'b1;
  assign CLBLM_R_X41Y92_SLICE_X66Y92_D6 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_A1 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_A2 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_A3 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_A4 = BRAM_L_X44Y95_RAMB18_X2Y38_DO9;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_A5 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_A6 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_AX = BRAM_L_X44Y95_RAMB18_X2Y38_DO7;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_B1 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_B2 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_B3 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_B4 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_B5 = BRAM_L_X44Y95_RAMB18_X2Y38_DOP0;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_B6 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_BX = BRAM_L_X44Y95_RAMB18_X2Y38_DO2;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_C1 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_C2 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_C3 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_C4 = BRAM_L_X44Y95_RAMB18_X2Y38_DO10;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_C5 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_C6 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_CE = CLBLL_L_X42Y97_SLICE_X69Y97_CO6;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_CX = BRAM_L_X44Y95_RAMB18_X2Y38_DO4;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_D1 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_D2 = BRAM_L_X44Y95_RAMB18_X2Y38_DO5;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_D3 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_D4 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_D5 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_D6 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X68Y111_DX = CLBLL_L_X42Y94_SLICE_X68Y94_BQ;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_A1 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_A2 = CLBLL_L_X42Y111_SLICE_X68Y111_BQ;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_A3 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_A4 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_A5 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_A6 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_AX = CLBLL_L_X42Y111_SLICE_X68Y111_A5Q;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_B1 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_B2 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_B3 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_B4 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_B5 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_B6 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_BX = CLBLL_L_X42Y98_SLICE_X69Y98_BQ;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_C1 = CLBLM_R_X41Y101_SLICE_X67Y101_DO6;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_C2 = CLBLM_R_X41Y106_SLICE_X67Y106_BO5;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_C3 = CLBLL_L_X42Y105_SLICE_X69Y105_BO5;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_C4 = CLBLM_R_X41Y101_SLICE_X67Y101_D5Q;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_C5 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_C6 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_CE = CLBLM_R_X41Y114_SLICE_X66Y114_DO6;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_D4 = CLBLM_R_X41Y101_SLICE_X67Y101_DQ;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_D1 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_D2 = CLBLL_L_X42Y111_SLICE_X68Y111_CQ;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_D3 = 1'b1;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_D5 = CLBLM_R_X41Y106_SLICE_X67Y106_BO6;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_D4 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_D5 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_D6 = 1'b1;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_D6 = 1'b1;
  assign CLBLL_L_X42Y111_SLICE_X69Y111_DX = CLBLL_L_X42Y111_SLICE_X68Y111_AQ;
  assign CLBLL_L_X42Y104_SLICE_X68Y104_DX = CLBLL_L_X42Y108_SLICE_X69Y108_CO5;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_A1 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_A2 = CLBLM_R_X41Y93_SLICE_X67Y93_AQ;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_A3 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_A4 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_A5 = CLBLM_R_X41Y95_SLICE_X67Y95_A_XOR;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_A6 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_AX = 1'b0;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_B1 = CLBLM_R_X41Y95_SLICE_X67Y95_C_XOR;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_B2 = CLBLM_R_X41Y93_SLICE_X67Y93_BQ;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_B3 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_B4 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_B5 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_B6 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_BX = 1'b0;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_C1 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_C2 = CLBLM_R_X41Y93_SLICE_X67Y93_CQ;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_C3 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_C4 = CLBLM_R_X41Y95_SLICE_X67Y95_D_XOR;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_C5 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_C6 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_CE = CLBLL_L_X42Y90_SLICE_X69Y90_CQ;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_CIN = CLBLM_R_X41Y92_SLICE_X67Y92_COUT;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_CX = 1'b0;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_D1 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_D2 = CLBLM_R_X41Y95_SLICE_X67Y95_B_XOR;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_D3 = CLBLM_R_X41Y93_SLICE_X67Y93_DQ;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_D4 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_D5 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_D6 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_DX = 1'b0;
  assign CLBLM_R_X41Y93_SLICE_X67Y93_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_A1 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_A2 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_A3 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_A4 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_A5 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_A6 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_B1 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_B2 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_B3 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_B4 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_B5 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_B6 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_C1 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_C2 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_C3 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_C4 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_C5 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_C6 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_D1 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_D2 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_D3 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_D4 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_D5 = 1'b1;
  assign CLBLM_R_X41Y93_SLICE_X66Y93_D6 = 1'b1;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_A1 = 1'b1;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_A2 = 1'b1;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_A4 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_C4 = 1'b1;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_A5 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_C5 = 1'b1;
  assign CLBLM_R_X3Y59_SLICE_X2Y59_C6 = 1'b1;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_AX = 1'b0;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_A1 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_A2 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_A3 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_A4 = CLBLL_L_X42Y91_SLICE_X68Y91_CQ;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_B1 = CLBLM_R_X41Y108_SLICE_X67Y108_BO6;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_A5 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_A6 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_AX = CLBLL_L_X42Y91_SLICE_X68Y91_AQ;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_B2 = CLBLL_L_X42Y104_SLICE_X69Y104_A_XOR;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_B1 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_B2 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_B3 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_B4 = 1'b1;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_B3 = CLBLL_L_X42Y103_SLICE_X68Y103_BQ;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_B5 = CLBLL_L_X42Y91_SLICE_X68Y91_BQ;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_B6 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_BX = CLBLL_L_X42Y90_SLICE_X68Y90_AQ;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_B4 = CLBLL_L_X42Y110_SLICE_X68Y110_BO5;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_C1 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_C2 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_C3 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_C4 = CLBLL_L_X42Y91_SLICE_X68Y91_DQ;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_B5 = 1'b0;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_C5 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_C6 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_CE = CLBLL_L_X42Y97_SLICE_X69Y97_CO6;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_B6 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_CX = CLBLL_L_X42Y90_SLICE_X68Y90_BQ;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_D1 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_D2 = CLBLL_L_X42Y90_SLICE_X68Y90_DQ;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_D3 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_D4 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_D5 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_D6 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X68Y112_DX = CLBLL_L_X42Y113_SLICE_X68Y113_D5Q;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_BX = 1'b0;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_C1 = CLBLL_L_X42Y103_SLICE_X69Y103_D_XOR;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR7 = CLBLL_L_X42Y90_SLICE_X68Y90_AQ;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_C2 = CLBLM_R_X41Y108_SLICE_X67Y108_BO6;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR8 = CLBLL_L_X42Y91_SLICE_X68Y91_AQ;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_C3 = 1'b0;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_C4 = CLBLL_L_X42Y110_SLICE_X68Y110_BO5;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_A1 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_A2 = CLBLL_L_X42Y71_SLICE_X68Y71_BQ;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_A3 = CLBLL_L_X42Y112_SLICE_X69Y112_BQ;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_A4 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_C5 = CLBLL_L_X42Y103_SLICE_X68Y103_CQ;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_A5 = CLBLL_L_X42Y112_SLICE_X69Y112_C5Q;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_A6 = CLBLL_L_X42Y43_SLICE_X68Y43_D_XOR;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR11 = CLBLL_L_X42Y91_SLICE_X68Y91_DQ;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_C6 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_B1 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_B2 = CLBLL_L_X42Y112_SLICE_X69Y112_DQ;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_B3 = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_ADDRARDADDR12 = CLBLL_L_X42Y92_SLICE_X69Y92_C5Q;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_CE = CLBLL_L_X42Y97_SLICE_X68Y97_CO6;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_B4 = CLBLL_L_X42Y112_SLICE_X69Y112_DO5;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_B5 = CLBLL_L_X42Y71_SLICE_X68Y71_BQ;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_B6 = 1'b1;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_CIN = CLBLL_L_X42Y103_SLICE_X69Y103_COUT;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_BX = CLBLL_L_X42Y112_SLICE_X69Y112_AO6;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_C1 = CLBLL_L_X42Y43_SLICE_X68Y43_D_XOR;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_C2 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_C3 = CLBLL_L_X42Y112_SLICE_X69Y112_DQ;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_C4 = CLBLL_L_X42Y112_SLICE_X69Y112_C5Q;
  assign CLBLL_L_X42Y104_SLICE_X69Y104_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_C5 = CLBLL_L_X42Y71_SLICE_X68Y71_BQ;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_C6 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_CLK = CLK_HROW_TOP_R_X78Y130_BUFHCE_X1Y34_O;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_D1 = CLBLL_L_X42Y94_SLICE_X69Y94_CQ;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_D2 = CLBLL_L_X42Y112_SLICE_X69Y112_BQ;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_D3 = CLBLL_L_X42Y71_SLICE_X68Y71_BQ;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_D4 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_D5 = CLBLL_L_X42Y110_SLICE_X69Y110_BQ;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_D6 = 1'b1;
  assign CLBLL_L_X42Y112_SLICE_X69Y112_DX = CLBLL_L_X42Y112_SLICE_X69Y112_BO5;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_A1 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_A2 = CLBLM_R_X41Y94_SLICE_X67Y94_CQ;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_A3 = CLBLM_R_X41Y94_SLICE_X67Y94_D_XOR;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_A4 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_A5 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_A6 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_AX = 1'b0;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_B1 = CLBLM_R_X41Y92_SLICE_X67Y92_D_XOR;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_B2 = CLBLM_R_X41Y94_SLICE_X67Y94_BQ;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_B3 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_B4 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_B5 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_B6 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_BX = 1'b0;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_C1 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_C2 = CLBLM_R_X41Y94_SLICE_X67Y94_DQ;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_C3 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_C4 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_C5 = CLBLM_R_X41Y94_SLICE_X67Y94_A_XOR;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_C6 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_CE = CLBLL_L_X42Y90_SLICE_X69Y90_CQ;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_CIN = CLBLM_R_X41Y93_SLICE_X67Y93_COUT;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_CLK = CLK_HROW_BOT_R_X78Y78_BUFHCE_X1Y20_O;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_CX = 1'b0;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_D1 = CLBLM_R_X41Y94_SLICE_X67Y94_C_XOR;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_D2 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_D3 = CLBLM_R_X41Y94_SLICE_X67Y94_AQ;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_D4 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_D5 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_D6 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_DX = 1'b0;
  assign CLBLM_R_X41Y94_SLICE_X67Y94_SR = CLBLL_L_X42Y96_SLICE_X69Y96_BO6;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_A1 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_A2 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_A3 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_A4 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_A5 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_A6 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_B1 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_B2 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_B3 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_B4 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_B5 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_B6 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_C1 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_C2 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_C3 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_C4 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_C5 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_C6 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_D1 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_D2 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_D3 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_D4 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_D5 = 1'b1;
  assign CLBLM_R_X41Y94_SLICE_X66Y94_D6 = 1'b1;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI14 = 1'b0;
  assign BRAM_L_X44Y95_RAMB18_X2Y38_DIADI15 = 1'b0;
endmodule
