// Copyright (C) 2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC

module top(
  input i_ce,
  input i_clk,
  input i_clkb,
  input i_rst,
  input [11:0] io,
  output o_q1,
  output o_q2
  );
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_A;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_A1;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_A2;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_A3;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_A4;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_A5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_A6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_AO5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_AO6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_A_CY;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_A_XOR;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_B;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_B1;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_B2;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_B3;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_B4;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_B5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_B6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_BO5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_BO6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_B_CY;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_B_XOR;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_C;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_C1;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_C2;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_C3;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_C4;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_C5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_C6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_CO5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_CO6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_C_CY;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_C_XOR;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_D;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_D1;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_D2;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_D3;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_D4;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_D5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_D6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_DO5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_DO6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_D_CY;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X0Y42_D_XOR;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_A;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_A1;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_A2;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_A3;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_A4;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_A5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_A6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_AMUX;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_AO5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_AO6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_A_CY;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_A_XOR;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_B;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_B1;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_B2;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_B3;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_B4;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_B5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_B6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_BMUX;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_BO5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_BO6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_B_CY;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_B_XOR;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_C;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_C1;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_C2;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_C3;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_C4;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_C5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_C6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_CMUX;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_CO5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_CO6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_C_CY;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_C_XOR;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_D;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_D1;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_D2;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_D3;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_D4;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_D5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_D6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_DO5;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_DO6;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_D_CY;
  wire [0:0] CLBLL_L_X2Y42_SLICE_X1Y42_D_XOR;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_A;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_A1;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_A2;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_A3;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_A4;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_A5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_A6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_AMUX;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_AO5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_AO6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_A_CY;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_A_XOR;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_B;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_B1;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_B2;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_B3;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_B4;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_B5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_B6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_BMUX;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_BO5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_BO6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_B_CY;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_B_XOR;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_C;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_C1;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_C2;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_C3;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_C4;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_C5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_C6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_CMUX;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_CO5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_CO6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_C_CY;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_C_XOR;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_D;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_D1;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_D2;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_D3;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_D4;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_D5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_D6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_DO5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_DO6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_D_CY;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X0Y43_D_XOR;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_A;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_A1;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_A2;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_A3;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_A4;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_A5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_A6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_AO5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_AO6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_A_CY;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_A_XOR;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_B;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_B1;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_B2;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_B3;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_B4;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_B5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_B6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_BO5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_BO6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_B_CY;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_B_XOR;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_C;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_C1;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_C2;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_C3;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_C4;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_C5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_C6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_CO5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_CO6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_C_CY;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_C_XOR;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_D;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_D1;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_D2;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_D3;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_D4;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_D5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_D6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_DO5;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_DO6;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_D_CY;
  wire [0:0] CLBLL_L_X2Y43_SLICE_X1Y43_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S1;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_CE;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_I;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_CE;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_I;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  wire [0:0] LIOB33_X0Y33_IOB_X0Y34_I;
  wire [0:0] LIOB33_X0Y35_IOB_X0Y35_I;
  wire [0:0] LIOB33_X0Y35_IOB_X0Y36_I;
  wire [0:0] LIOB33_X0Y37_IOB_X0Y37_I;
  wire [0:0] LIOB33_X0Y37_IOB_X0Y38_I;
  wire [0:0] LIOB33_X0Y39_IOB_X0Y39_I;
  wire [0:0] LIOB33_X0Y39_IOB_X0Y40_I;
  wire [0:0] LIOB33_X0Y41_IOB_X0Y41_I;
  wire [0:0] LIOB33_X0Y41_IOB_X0Y42_I;
  wire [0:0] LIOB33_X0Y43_IOB_X0Y43_I;
  wire [0:0] LIOB33_X0Y45_IOB_X0Y45_I;
  wire [0:0] LIOB33_X0Y45_IOB_X0Y46_I;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_CE1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_CLK;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_CLKB;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q2;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_SR;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_CE1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_CLK;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_CLKB;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q2;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_SR;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_CE1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_CLK;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_CLKB;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q2;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_SR;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y34_CE1;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y34_CLK;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y34_CLKB;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y34_D;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y34_Q1;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y34_Q2;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y34_SR;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y35_CE1;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y35_CLK;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y35_CLKB;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y35_D;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y35_Q1;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y35_Q2;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y35_SR;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y36_CE1;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y36_CLK;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y36_CLKB;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y36_D;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y36_Q1;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y36_Q2;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y36_SR;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y39_CE1;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y39_CLK;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y39_CLKB;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y39_D;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y39_Q1;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y39_Q2;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y39_SR;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y40_CE1;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y40_CLK;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y40_CLKB;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y40_D;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y40_Q1;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y40_Q2;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y40_SR;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y41_CE1;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y41_CLK;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y41_CLKB;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y41_D;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y41_Q1;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y41_Q2;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y41_SR;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y42_CE1;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y42_CLK;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y42_CLKB;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y42_D;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y42_Q1;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y42_Q2;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y42_SR;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y45_CE1;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y45_CLK;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y45_CLKB;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y45_D;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y45_Q1;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y45_Q2;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y45_SR;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y46_CE1;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y46_CLK;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y46_CLKB;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y46_D;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y46_Q1;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y46_Q2;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y46_SR;
  wire [0:0] RIOB33_X43Y23_IOB_X1Y24_I;
  wire [0:0] RIOB33_X43Y25_IOB_X1Y26_I;
  wire [0:0] RIOB33_X43Y43_IOB_X1Y43_O;
  wire [0:0] RIOB33_X43Y43_IOB_X1Y44_O;
  wire [0:0] RIOB33_X43Y45_IOB_X1Y45_I;
  wire [0:0] RIOB33_X43Y45_IOB_X1Y46_I;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_D1;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_OQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_T1;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_TQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_D1;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_OQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_T1;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_TQ;
  wire [0:0] RIOI3_X43Y23_ILOGIC_X1Y24_D;
  wire [0:0] RIOI3_X43Y23_ILOGIC_X1Y24_O;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_D;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_O;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y45_D;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y45_O;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y46_D;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y46_O;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y42_SLICE_X0Y42_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y42_SLICE_X0Y42_DO5),
.O6(CLBLL_L_X2Y42_SLICE_X0Y42_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y42_SLICE_X0Y42_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y42_SLICE_X0Y42_CO5),
.O6(CLBLL_L_X2Y42_SLICE_X0Y42_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y42_SLICE_X0Y42_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y42_SLICE_X0Y42_BO5),
.O6(CLBLL_L_X2Y42_SLICE_X0Y42_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y42_SLICE_X0Y42_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y42_SLICE_X0Y42_AO5),
.O6(CLBLL_L_X2Y42_SLICE_X0Y42_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y42_SLICE_X1Y42_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y42_SLICE_X1Y42_DO5),
.O6(CLBLL_L_X2Y42_SLICE_X1Y42_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010100000000)
  ) CLBLL_L_X2Y42_SLICE_X1Y42_CLUT (
.I0(LIOI3_X0Y35_ILOGIC_X0Y36_Q1),
.I1(LIOI3_X0Y33_ILOGIC_X0Y34_Q1),
.I2(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q1),
.I3(1'b1),
.I4(LIOI3_X0Y35_ILOGIC_X0Y35_Q1),
.I5(1'b1),
.O5(CLBLL_L_X2Y42_SLICE_X1Y42_CO5),
.O6(CLBLL_L_X2Y42_SLICE_X1Y42_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000500000000)
  ) CLBLL_L_X2Y42_SLICE_X1Y42_BLUT (
.I0(LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q1),
.I1(1'b1),
.I2(LIOI3_X0Y45_ILOGIC_X0Y45_Q1),
.I3(LIOI3_X0Y41_ILOGIC_X0Y42_Q1),
.I4(LIOI3_X0Y45_ILOGIC_X0Y46_Q1),
.I5(1'b1),
.O5(CLBLL_L_X2Y42_SLICE_X1Y42_BO5),
.O6(CLBLL_L_X2Y42_SLICE_X1Y42_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdffffffff)
  ) CLBLL_L_X2Y42_SLICE_X1Y42_ALUT (
.I0(CLBLL_L_X2Y42_SLICE_X1Y42_BO6),
.I1(LIOI3_X0Y39_ILOGIC_X0Y39_Q1),
.I2(LIOI3_X0Y41_ILOGIC_X0Y41_Q1),
.I3(LIOI3_X0Y39_ILOGIC_X0Y40_Q1),
.I4(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q1),
.I5(CLBLL_L_X2Y42_SLICE_X1Y42_CO6),
.O5(CLBLL_L_X2Y42_SLICE_X1Y42_AO5),
.O6(CLBLL_L_X2Y42_SLICE_X1Y42_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y43_SLICE_X0Y43_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y43_SLICE_X0Y43_DO5),
.O6(CLBLL_L_X2Y43_SLICE_X0Y43_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010100000000)
  ) CLBLL_L_X2Y43_SLICE_X0Y43_CLUT (
.I0(LIOI3_X0Y35_ILOGIC_X0Y36_Q2),
.I1(LIOI3_X0Y33_ILOGIC_X0Y34_Q2),
.I2(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q2),
.I3(1'b1),
.I4(LIOI3_X0Y35_ILOGIC_X0Y35_Q2),
.I5(1'b1),
.O5(CLBLL_L_X2Y43_SLICE_X0Y43_CO5),
.O6(CLBLL_L_X2Y43_SLICE_X0Y43_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000500000000)
  ) CLBLL_L_X2Y43_SLICE_X0Y43_BLUT (
.I0(LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q2),
.I1(1'b1),
.I2(LIOI3_X0Y45_ILOGIC_X0Y45_Q2),
.I3(LIOI3_X0Y41_ILOGIC_X0Y42_Q2),
.I4(LIOI3_X0Y45_ILOGIC_X0Y46_Q2),
.I5(1'b1),
.O5(CLBLL_L_X2Y43_SLICE_X0Y43_BO5),
.O6(CLBLL_L_X2Y43_SLICE_X0Y43_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdffffffff)
  ) CLBLL_L_X2Y43_SLICE_X0Y43_ALUT (
.I0(CLBLL_L_X2Y43_SLICE_X0Y43_BO6),
.I1(LIOI3_X0Y39_ILOGIC_X0Y39_Q2),
.I2(LIOI3_X0Y41_ILOGIC_X0Y41_Q2),
.I3(LIOI3_X0Y39_ILOGIC_X0Y40_Q2),
.I4(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q2),
.I5(CLBLL_L_X2Y43_SLICE_X0Y43_CO6),
.O5(CLBLL_L_X2Y43_SLICE_X0Y43_AO5),
.O6(CLBLL_L_X2Y43_SLICE_X0Y43_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y43_SLICE_X1Y43_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y43_SLICE_X1Y43_DO5),
.O6(CLBLL_L_X2Y43_SLICE_X1Y43_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y43_SLICE_X1Y43_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y43_SLICE_X1Y43_CO5),
.O6(CLBLL_L_X2Y43_SLICE_X1Y43_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y43_SLICE_X1Y43_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y43_SLICE_X1Y43_BO5),
.O6(CLBLL_L_X2Y43_SLICE_X1Y43_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y43_SLICE_X1Y43_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y43_SLICE_X1Y43_AO5),
.O6(CLBLL_L_X2Y43_SLICE_X1Y43_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X43Y25_IOB_X1Y26_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X43Y23_IOB_X1Y24_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O),
.O(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y33_IOB_X0Y34_IBUF (
.I(io[11]),
.O(LIOB33_X0Y33_IOB_X0Y34_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y35_IOB_X0Y35_IBUF (
.I(io[10]),
.O(LIOB33_X0Y35_IOB_X0Y35_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y35_IOB_X0Y36_IBUF (
.I(io[9]),
.O(LIOB33_X0Y35_IOB_X0Y36_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y37_IOB_X0Y37_IBUF (
.I(io[8]),
.O(LIOB33_X0Y37_IOB_X0Y37_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y37_IOB_X0Y38_IBUF (
.I(io[7]),
.O(LIOB33_X0Y37_IOB_X0Y38_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y39_IOB_X0Y39_IBUF (
.I(io[6]),
.O(LIOB33_X0Y39_IOB_X0Y39_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y39_IOB_X0Y40_IBUF (
.I(io[5]),
.O(LIOB33_X0Y39_IOB_X0Y40_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y41_IOB_X0Y41_IBUF (
.I(io[4]),
.O(LIOB33_X0Y41_IOB_X0Y41_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y41_IOB_X0Y42_IBUF (
.I(io[3]),
.O(LIOB33_X0Y41_IOB_X0Y42_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y43_IOB_X0Y43_IBUF (
.I(io[2]),
.O(LIOB33_X0Y43_IOB_X0Y43_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y45_IOB_X0Y45_IBUF (
.I(io[1]),
.O(LIOB33_X0Y45_IOB_X0Y45_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y45_IOB_X0Y46_IBUF (
.I(io[0]),
.O(LIOB33_X0Y45_IOB_X0Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b1),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y33_ILOGIC_X0Y34_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y33_IOB_X0Y34_I),
.Q1(LIOI3_X0Y33_ILOGIC_X0Y34_Q1),
.Q2(LIOI3_X0Y33_ILOGIC_X0Y34_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y35_ILOGIC_X0Y36_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y35_IOB_X0Y36_I),
.Q1(LIOI3_X0Y35_ILOGIC_X0Y36_Q1),
.Q2(LIOI3_X0Y35_ILOGIC_X0Y36_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y35_ILOGIC_X0Y35_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y35_IOB_X0Y35_I),
.Q1(LIOI3_X0Y35_ILOGIC_X0Y35_Q1),
.Q2(LIOI3_X0Y35_ILOGIC_X0Y35_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y39_ILOGIC_X0Y40_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y39_IOB_X0Y40_I),
.Q1(LIOI3_X0Y39_ILOGIC_X0Y40_Q1),
.Q2(LIOI3_X0Y39_ILOGIC_X0Y40_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y39_ILOGIC_X0Y39_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y39_IOB_X0Y39_I),
.Q1(LIOI3_X0Y39_ILOGIC_X0Y39_Q1),
.Q2(LIOI3_X0Y39_ILOGIC_X0Y39_Q2),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE_PIPELINED"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y41_ILOGIC_X0Y42_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y41_IOB_X0Y42_I),
.Q1(LIOI3_X0Y41_ILOGIC_X0Y42_Q1),
.Q2(LIOI3_X0Y41_ILOGIC_X0Y42_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y41_ILOGIC_X0Y41_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y41_IOB_X0Y41_I),
.Q1(LIOI3_X0Y41_ILOGIC_X0Y41_Q1),
.Q2(LIOI3_X0Y41_ILOGIC_X0Y41_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y45_ILOGIC_X0Y46_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y45_IOB_X0Y46_I),
.Q1(LIOI3_X0Y45_ILOGIC_X0Y46_Q1),
.Q2(LIOI3_X0Y45_ILOGIC_X0Y46_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y45_ILOGIC_X0Y45_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y45_IOB_X0Y45_I),
.Q1(LIOI3_X0Y45_ILOGIC_X0Y45_Q1),
.Q2(LIOI3_X0Y45_ILOGIC_X0Y45_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y43_IOB_X0Y43_I),
.Q1(LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q1),
.Q2(LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y37_IOB_X0Y38_I),
.Q1(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q1),
.Q2(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q2),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y37_IOB_X0Y37_I),
.Q1(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q1),
.Q2(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y23_IOB_X1Y24_IBUF (
.I(i_clkb),
.O(RIOB33_X43Y23_IOB_X1Y24_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y25_IOB_X1Y26_IBUF (
.I(i_clk),
.O(RIOB33_X43Y25_IOB_X1Y26_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y43_IOB_X1Y43_OBUF (
.I(CLBLL_L_X2Y43_SLICE_X0Y43_AO6),
.O(o_q2)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y43_IOB_X1Y44_OBUF (
.I(CLBLL_L_X2Y42_SLICE_X1Y42_AO6),
.O(o_q1)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y45_IOB_X1Y45_IBUF (
.I(i_ce),
.O(RIOB33_X43Y45_IOB_X1Y45_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y45_IOB_X1Y46_IBUF (
.I(i_rst),
.O(RIOB33_X43Y45_IOB_X1Y46_I)
  );
  assign CLBLL_L_X2Y42_SLICE_X0Y42_A = CLBLL_L_X2Y42_SLICE_X0Y42_AO6;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_B = CLBLL_L_X2Y42_SLICE_X0Y42_BO6;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_C = CLBLL_L_X2Y42_SLICE_X0Y42_CO6;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_D = CLBLL_L_X2Y42_SLICE_X0Y42_DO6;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_A = CLBLL_L_X2Y42_SLICE_X1Y42_AO6;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_B = CLBLL_L_X2Y42_SLICE_X1Y42_BO6;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_C = CLBLL_L_X2Y42_SLICE_X1Y42_CO6;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_D = CLBLL_L_X2Y42_SLICE_X1Y42_DO6;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_AMUX = CLBLL_L_X2Y42_SLICE_X1Y42_AO6;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_BMUX = CLBLL_L_X2Y42_SLICE_X1Y42_BO6;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_CMUX = CLBLL_L_X2Y42_SLICE_X1Y42_CO6;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_A = CLBLL_L_X2Y43_SLICE_X0Y43_AO6;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_B = CLBLL_L_X2Y43_SLICE_X0Y43_BO6;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_C = CLBLL_L_X2Y43_SLICE_X0Y43_CO6;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_D = CLBLL_L_X2Y43_SLICE_X0Y43_DO6;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_AMUX = CLBLL_L_X2Y43_SLICE_X0Y43_AO6;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_BMUX = CLBLL_L_X2Y43_SLICE_X0Y43_BO6;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_CMUX = CLBLL_L_X2Y43_SLICE_X0Y43_CO6;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_A = CLBLL_L_X2Y43_SLICE_X1Y43_AO6;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_B = CLBLL_L_X2Y43_SLICE_X1Y43_BO6;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_C = CLBLL_L_X2Y43_SLICE_X1Y43_CO6;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_D = CLBLL_L_X2Y43_SLICE_X1Y43_DO6;
  assign RIOI3_X43Y23_ILOGIC_X1Y24_O = RIOB33_X43Y23_IOB_X1Y24_I;
  assign RIOI3_X43Y25_ILOGIC_X1Y26_O = RIOB33_X43Y25_IOB_X1Y26_I;
  assign RIOI3_X43Y45_ILOGIC_X1Y46_O = RIOB33_X43Y45_IOB_X1Y46_I;
  assign RIOI3_X43Y45_ILOGIC_X1Y45_O = RIOB33_X43Y45_IOB_X1Y45_I;
  assign RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_OQ = CLBLL_L_X2Y42_SLICE_X1Y42_AO6;
  assign RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_OQ = CLBLL_L_X2Y43_SLICE_X0Y43_AO6;
  assign RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_D1 = CLBLL_L_X2Y42_SLICE_X1Y42_AO6;
  assign LIOI3_X0Y39_ILOGIC_X0Y40_D = LIOB33_X0Y39_IOB_X0Y40_I;
  assign LIOI3_X0Y39_ILOGIC_X0Y39_D = LIOB33_X0Y39_IOB_X0Y39_I;
  assign LIOI3_X0Y39_ILOGIC_X0Y40_SR = 1'b0;
  assign LIOI3_X0Y39_ILOGIC_X0Y39_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y39_ILOGIC_X0Y39_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y39_ILOGIC_X0Y39_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_T1 = 1'b1;
  assign RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_D1 = CLBLL_L_X2Y43_SLICE_X0Y43_AO6;
  assign LIOI3_X0Y39_ILOGIC_X0Y39_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y33_ILOGIC_X0Y34_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_T1 = 1'b1;
  assign LIOI3_X0Y33_ILOGIC_X0Y34_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y33_ILOGIC_X0Y34_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign LIOI3_X0Y33_ILOGIC_X0Y34_D = LIOB33_X0Y33_IOB_X0Y34_I;
  assign RIOI3_X43Y23_ILOGIC_X1Y24_D = RIOB33_X43Y23_IOB_X1Y24_I;
  assign LIOI3_X0Y33_ILOGIC_X0Y34_SR = 1'b0;
  assign LIOI3_X0Y41_ILOGIC_X0Y41_SR = 1'b0;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_A1 = CLBLL_L_X2Y43_SLICE_X0Y43_BO6;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_A2 = LIOI3_X0Y39_ILOGIC_X0Y39_Q2;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_A3 = LIOI3_X0Y41_ILOGIC_X0Y41_Q2;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_A4 = LIOI3_X0Y39_ILOGIC_X0Y40_Q2;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_A5 = LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q2;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_A6 = CLBLL_L_X2Y43_SLICE_X0Y43_CO6;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_B1 = LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q2;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_B2 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_B3 = LIOI3_X0Y45_ILOGIC_X0Y45_Q2;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_B4 = LIOI3_X0Y41_ILOGIC_X0Y42_Q2;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_B5 = LIOI3_X0Y45_ILOGIC_X0Y46_Q2;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_B6 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_C1 = LIOI3_X0Y35_ILOGIC_X0Y36_Q2;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_C2 = LIOI3_X0Y33_ILOGIC_X0Y34_Q2;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_C3 = LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q2;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_C4 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_C5 = LIOI3_X0Y35_ILOGIC_X0Y35_Q2;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_C6 = 1'b1;
  assign LIOI3_X0Y35_ILOGIC_X0Y36_SR = 1'b0;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_D1 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_D2 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_D3 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_D4 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_D5 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X0Y43_D6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_D = LIOB33_X0Y37_IOB_X0Y38_I;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_D = LIOB33_X0Y37_IOB_X0Y37_I;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign LIOI3_X0Y41_ILOGIC_X0Y42_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y41_ILOGIC_X0Y42_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y41_ILOGIC_X0Y42_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_A1 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_A2 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_A3 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_A4 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_A5 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_A6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_SR = 1'b0;
  assign LIOI3_X0Y41_ILOGIC_X0Y42_D = LIOB33_X0Y41_IOB_X0Y42_I;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_B1 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_B2 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_B3 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_B4 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_B5 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_B6 = 1'b1;
  assign LIOI3_X0Y41_ILOGIC_X0Y42_SR = 1'b0;
  assign LIOI3_X0Y41_ILOGIC_X0Y41_D = LIOB33_X0Y41_IOB_X0Y41_I;
  assign LIOI3_X0Y41_ILOGIC_X0Y41_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_C1 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_C2 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_C3 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_C4 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_C5 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_C6 = 1'b1;
  assign LIOI3_X0Y41_ILOGIC_X0Y41_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y41_ILOGIC_X0Y41_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_D1 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_D2 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_D3 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_D4 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_D5 = 1'b1;
  assign CLBLL_L_X2Y43_SLICE_X1Y43_D6 = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_CE = 1'b1;
  assign LIOI3_X0Y35_ILOGIC_X0Y36_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_CE = 1'b1;
  assign LIOI3_X0Y35_ILOGIC_X0Y36_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y35_ILOGIC_X0Y36_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign LIOI3_X0Y35_ILOGIC_X0Y36_D = LIOB33_X0Y35_IOB_X0Y36_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign LIOI3_X0Y35_ILOGIC_X0Y35_D = LIOB33_X0Y35_IOB_X0Y35_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S1 = 1'b1;
  assign LIOI3_X0Y35_ILOGIC_X0Y35_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y35_ILOGIC_X0Y35_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y35_ILOGIC_X0Y35_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign LIOI3_X0Y35_ILOGIC_X0Y35_SR = 1'b0;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_A1 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_A2 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_A3 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_A4 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_A5 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_A6 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_B1 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_B2 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_B3 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_B4 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_B5 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_B6 = 1'b1;
  assign RIOI3_X43Y45_ILOGIC_X1Y46_D = RIOB33_X43Y45_IOB_X1Y46_I;
  assign RIOI3_X43Y45_ILOGIC_X1Y45_D = RIOB33_X43Y45_IOB_X1Y45_I;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_C1 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_C2 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_C3 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_C4 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_C5 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_C6 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_D1 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_D2 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_D3 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_D4 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_D5 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X0Y42_D6 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0 = RIOB33_X43Y25_IOB_X1Y26_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_A1 = CLBLL_L_X2Y42_SLICE_X1Y42_BO6;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I0 = RIOB33_X43Y23_IOB_X1Y24_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I1 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_A2 = LIOI3_X0Y39_ILOGIC_X0Y39_Q1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_A3 = LIOI3_X0Y41_ILOGIC_X0Y41_Q1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_A4 = LIOI3_X0Y39_ILOGIC_X0Y40_Q1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_A5 = LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_A6 = CLBLL_L_X2Y42_SLICE_X1Y42_CO6;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_B1 = LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_B2 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_B3 = LIOI3_X0Y45_ILOGIC_X0Y45_Q1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_B4 = LIOI3_X0Y41_ILOGIC_X0Y42_Q1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_B5 = LIOI3_X0Y45_ILOGIC_X0Y46_Q1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_B6 = 1'b1;
  assign RIOI3_X43Y25_ILOGIC_X1Y26_D = RIOB33_X43Y25_IOB_X1Y26_I;
  assign LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_D = LIOB33_X0Y43_IOB_X0Y43_I;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_C1 = LIOI3_X0Y35_ILOGIC_X0Y36_Q1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_C2 = LIOI3_X0Y33_ILOGIC_X0Y34_Q1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_C3 = LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_C4 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_C5 = LIOI3_X0Y35_ILOGIC_X0Y35_Q1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_C6 = 1'b1;
  assign LIOI3_X0Y45_ILOGIC_X0Y46_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y45_ILOGIC_X0Y46_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y45_ILOGIC_X0Y46_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_D1 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_D2 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_D3 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_D4 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_D5 = 1'b1;
  assign CLBLL_L_X2Y42_SLICE_X1Y42_D6 = 1'b1;
  assign LIOI3_X0Y45_ILOGIC_X0Y46_D = LIOB33_X0Y45_IOB_X0Y46_I;
  assign LIOI3_X0Y45_ILOGIC_X0Y45_D = LIOB33_X0Y45_IOB_X0Y45_I;
  assign LIOI3_X0Y45_ILOGIC_X0Y46_SR = 1'b0;
  assign LIOI3_X0Y45_ILOGIC_X0Y45_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_SR = 1'b0;
  assign LIOI3_X0Y45_ILOGIC_X0Y45_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y45_ILOGIC_X0Y45_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign RIOB33_X43Y43_IOB_X1Y43_O = CLBLL_L_X2Y43_SLICE_X0Y43_AO6;
  assign RIOB33_X43Y43_IOB_X1Y44_O = CLBLL_L_X2Y42_SLICE_X1Y42_AO6;
  assign LIOI3_X0Y45_ILOGIC_X0Y45_SR = 1'b0;
  assign LIOI3_X0Y39_ILOGIC_X0Y40_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y39_ILOGIC_X0Y40_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y39_ILOGIC_X0Y40_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
endmodule
