module top(
  input clk,
  input jc4,
  input [7:0] sw,
  output jc2,
  output [7:0] led
  );
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_A;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_A1;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_A2;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_A3;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_A4;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_A5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_A6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_AMUX;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_AO5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_AO6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_A_CY;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_A_XOR;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_B;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_B1;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_B2;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_B3;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_B4;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_B5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_B6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_BO5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_BO6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_B_CY;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_B_XOR;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_C;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_C1;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_C2;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_C3;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_C4;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_C5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_C6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_CLK;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_CO5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_CO6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_C_CY;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_C_XOR;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_D;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_D1;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_D2;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_D3;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_D4;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_D5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_D6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_DO5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_DO6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_DQ;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_DX;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_D_CY;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X36Y46_D_XOR;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_A;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_A1;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_A2;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_A3;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_A4;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_A5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_A6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_AO5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_AO6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_A_CY;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_A_XOR;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_B;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_B1;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_B2;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_B3;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_B4;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_B5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_B6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_BO5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_BO6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_B_CY;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_B_XOR;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_C;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_C1;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_C2;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_C3;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_C4;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_C5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_C6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_CO5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_CO6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_C_CY;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_C_XOR;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_D;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_D1;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_D2;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_D3;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_D4;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_D5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_D6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_DO5;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_DO6;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_D_CY;
  wire [0:0] CLBLL_L_X24Y46_SLICE_X37Y46_D_XOR;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_A;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_A1;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_A2;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_A3;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_A4;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_A5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_A6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_AO5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_AO6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_A_CY;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_A_XOR;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_B;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_B1;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_B2;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_B3;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_B4;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_B5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_B6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_BO5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_BO6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_B_CY;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_B_XOR;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_C;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_C1;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_C2;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_C3;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_C4;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_C5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_C6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_CLK;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_CO5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_CO6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_C_CY;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_C_XOR;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_D;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_D1;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_D2;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_D3;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_D4;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_D5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_D6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_DO5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_DO6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_DQ;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_DX;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_D_CY;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X40Y9_D_XOR;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_A;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_A1;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_A2;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_A3;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_A4;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_A5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_A6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_AO5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_AO6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_A_CY;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_A_XOR;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_B;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_B1;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_B2;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_B3;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_B4;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_B5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_B6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_BO5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_BO6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_B_CY;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_B_XOR;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_C;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_C1;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_C2;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_C3;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_C4;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_C5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_C6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_CO5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_CO6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_C_CY;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_C_XOR;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_D;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_D1;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_D2;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_D3;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_D4;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_D5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_D6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_DO5;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_DO6;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_D_CY;
  wire [0:0] CLBLL_L_X26Y9_SLICE_X41Y9_D_XOR;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_A;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_A1;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_A2;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_A3;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_A4;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_A5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_A6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_AO5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_AO6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_A_CY;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_A_XOR;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_B;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_B1;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_B2;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_B3;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_B4;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_B5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_B6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_BO5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_BO6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_B_CY;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_B_XOR;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_C;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_C1;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_C2;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_C3;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_C4;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_C5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_C6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_CO5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_CO6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_C_CY;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_C_XOR;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_D;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_D1;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_D2;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_D3;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_D4;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_D5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_D6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_DO5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_DO6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_D_CY;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X14Y10_D_XOR;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_A;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_A1;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_A2;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_A3;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_A4;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_A5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_A6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_AMUX;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_AO5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_AO6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_AQ;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_AX;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_A_CY;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_A_XOR;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_B;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_B1;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_B2;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_B3;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_B4;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_B5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_B6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_BMUX;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_BO5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_BO6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_BQ;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_BX;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_B_CY;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_B_XOR;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_C;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_C1;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_C2;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_C3;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_C4;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_C5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_C6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_CIN;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_CLK;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_CO5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_CO6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_COUT;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_CQ;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_CX;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_C_CY;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_C_XOR;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_D;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_D1;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_D2;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_D3;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_D4;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_D5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_D6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_DO5;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_DO6;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_DQ;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_DX;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_D_CY;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_D_XOR;
  wire [0:0] CLBLM_R_X11Y10_SLICE_X15Y10_SR;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_A;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_A1;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_A2;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_A3;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_A4;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_A5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_A6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_AMUX;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_AO5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_AO6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_AQ;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_AX;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_A_CY;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_A_XOR;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_B;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_B1;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_B2;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_B3;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_B4;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_B5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_B6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_BMUX;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_BO5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_BO6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_BQ;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_BX;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_B_CY;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_B_XOR;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_C;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_C1;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_C2;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_C3;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_C4;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_C5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_C6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_CLK;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_CMUX;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_CO5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_CO6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_COUT;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_CQ;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_CX;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_C_CY;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_C_XOR;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_D;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_D1;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_D2;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_D3;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_D4;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_D5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_D6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_DMUX;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_DO5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_DO6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_DQ;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_DX;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_D_CY;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_D_XOR;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X14Y28_SR;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_A;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_A1;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_A2;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_A3;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_A4;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_A5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_A6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_AO5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_AO6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_A_CY;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_A_XOR;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_B;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_B1;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_B2;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_B3;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_B4;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_B5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_B6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_BO5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_BO6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_B_CY;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_B_XOR;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_C;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_C1;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_C2;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_C3;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_C4;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_C5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_C6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_CO5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_CO6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_C_CY;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_C_XOR;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_D;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_D1;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_D2;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_D3;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_D4;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_D5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_D6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_DO5;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_DO6;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_D_CY;
  wire [0:0] CLBLM_R_X11Y28_SLICE_X15Y28_D_XOR;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_A;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_A1;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_A2;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_A3;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_A4;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_A5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_A6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_AMUX;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_AO5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_AO6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_AQ;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_AX;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_A_CY;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_A_XOR;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_B;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_B1;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_B2;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_B3;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_B4;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_B5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_B6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_BMUX;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_BO5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_BO6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_BQ;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_BX;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_B_CY;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_B_XOR;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_C;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_C1;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_C2;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_C3;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_C4;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_C5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_C6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_CIN;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_CLK;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_CMUX;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_CO5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_CO6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_COUT;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_CQ;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_CX;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_C_CY;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_C_XOR;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_D;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_D1;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_D2;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_D3;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_D4;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_D5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_D6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_DMUX;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_DO5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_DO6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_DQ;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_DX;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_D_CY;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_D_XOR;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X14Y29_SR;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_A;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_A1;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_A2;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_A3;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_A4;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_A5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_A6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_AO5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_AO6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_A_CY;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_A_XOR;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_B;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_B1;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_B2;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_B3;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_B4;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_B5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_B6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_BO5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_BO6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_B_CY;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_B_XOR;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_C;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_C1;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_C2;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_C3;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_C4;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_C5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_C6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_CO5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_CO6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_C_CY;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_C_XOR;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_D;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_D1;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_D2;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_D3;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_D4;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_D5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_D6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_DO5;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_DO6;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_D_CY;
  wire [0:0] CLBLM_R_X11Y29_SLICE_X15Y29_D_XOR;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_A;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_A1;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_A2;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_A3;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_A4;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_A5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_A6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_AMUX;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_AO5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_AO6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_AQ;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_AX;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_A_CY;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_A_XOR;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_B;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_B1;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_B2;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_B3;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_B4;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_B5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_B6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_BMUX;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_BO5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_BO6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_BQ;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_BX;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_B_CY;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_B_XOR;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_C;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_C1;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_C2;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_C3;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_C4;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_C5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_C6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_CIN;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_CLK;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_CMUX;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_CO5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_CO6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_COUT;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_CQ;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_CX;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_C_CY;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_C_XOR;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_D;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_D1;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_D2;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_D3;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_D4;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_D5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_D6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_DMUX;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_DO5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_DO6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_DQ;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_DX;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_D_CY;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_D_XOR;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X14Y30_SR;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_A;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_A1;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_A2;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_A3;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_A4;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_A5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_A6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_AO5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_AO6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_A_CY;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_A_XOR;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_B;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_B1;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_B2;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_B3;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_B4;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_B5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_B6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_BO5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_BO6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_B_CY;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_B_XOR;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_C;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_C1;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_C2;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_C3;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_C4;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_C5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_C6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_CO5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_CO6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_C_CY;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_C_XOR;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_D;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_D1;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_D2;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_D3;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_D4;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_D5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_D6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_DO5;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_DO6;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_D_CY;
  wire [0:0] CLBLM_R_X11Y30_SLICE_X15Y30_D_XOR;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_A;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_A1;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_A2;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_A3;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_A4;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_A5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_A6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_AO5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_AO6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_AQ;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_AX;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_A_CY;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_A_XOR;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_B;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_B1;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_B2;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_B3;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_B4;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_B5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_B6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_BMUX;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_BO5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_BO6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_BQ;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_BX;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_B_CY;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_B_XOR;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_C;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_C1;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_C2;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_C3;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_C4;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_C5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_C6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_CIN;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_CLK;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_CMUX;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_CO5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_CO6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_COUT;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_CQ;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_CX;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_C_CY;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_C_XOR;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_D;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_D1;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_D2;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_D3;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_D4;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_D5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_D6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_DMUX;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_DO5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_DO6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_DQ;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_DX;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_D_CY;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_D_XOR;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X14Y31_SR;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_A;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_A1;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_A2;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_A3;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_A4;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_A5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_A6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_AO5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_AO6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_A_CY;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_A_XOR;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_B;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_B1;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_B2;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_B3;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_B4;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_B5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_B6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_BO5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_BO6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_B_CY;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_B_XOR;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_C;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_C1;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_C2;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_C3;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_C4;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_C5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_C6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_CO5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_CO6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_C_CY;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_C_XOR;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_D;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_D1;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_D2;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_D3;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_D4;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_D5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_D6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_DO5;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_DO6;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_D_CY;
  wire [0:0] CLBLM_R_X11Y31_SLICE_X15Y31_D_XOR;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_A;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_A1;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_A2;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_A3;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_A4;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_A5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_A6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_AO5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_AO6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_AQ;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_AX;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_A_CY;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_A_XOR;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_B;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_B1;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_B2;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_B3;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_B4;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_B5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_B6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_BMUX;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_BO5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_BO6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_BQ;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_BX;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_B_CY;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_B_XOR;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_C;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_C1;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_C2;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_C3;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_C4;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_C5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_C6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_CIN;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_CLK;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_CMUX;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_CO5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_CO6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_COUT;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_CQ;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_CX;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_C_CY;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_C_XOR;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_D;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_D1;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_D2;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_D3;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_D4;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_D5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_D6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_DMUX;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_DO5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_DO6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_DQ;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_DX;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_D_CY;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_D_XOR;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X14Y32_SR;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_A;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_A1;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_A2;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_A3;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_A4;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_A5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_A6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_AO5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_AO6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_A_CY;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_A_XOR;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_B;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_B1;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_B2;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_B3;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_B4;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_B5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_B6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_BO5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_BO6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_B_CY;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_B_XOR;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_C;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_C1;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_C2;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_C3;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_C4;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_C5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_C6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_CO5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_CO6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_C_CY;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_C_XOR;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_D;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_D1;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_D2;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_D3;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_D4;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_D5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_D6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_DO5;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_DO6;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_D_CY;
  wire [0:0] CLBLM_R_X11Y32_SLICE_X15Y32_D_XOR;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_A;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_A1;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_A2;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_A3;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_A4;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_A5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_A6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_AMUX;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_AO5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_AO6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_AQ;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_AX;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_A_CY;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_A_XOR;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_B;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_B1;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_B2;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_B3;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_B4;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_B5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_B6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_BMUX;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_BO5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_BO6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_BQ;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_BX;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_B_CY;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_B_XOR;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_C;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_C1;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_C2;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_C3;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_C4;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_C5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_C6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_CIN;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_CLK;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_CO5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_CO6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_COUT;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_CQ;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_CX;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_C_CY;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_C_XOR;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_D;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_D1;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_D2;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_D3;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_D4;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_D5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_D6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_DO5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_DO6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_DQ;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_DX;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_D_CY;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_D_XOR;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X14Y33_SR;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_A;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_A1;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_A2;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_A3;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_A4;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_A5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_A6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_AO5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_AO6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_A_CY;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_A_XOR;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_B;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_B1;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_B2;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_B3;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_B4;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_B5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_B6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_BO5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_BO6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_B_CY;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_B_XOR;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_C;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_C1;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_C2;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_C3;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_C4;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_C5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_C6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_CO5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_CO6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_C_CY;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_C_XOR;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_D;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_D1;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_D2;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_D3;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_D4;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_D5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_D6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_DO5;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_DO6;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_D_CY;
  wire [0:0] CLBLM_R_X11Y33_SLICE_X15Y33_D_XOR;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_A;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_A1;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_A2;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_A3;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_A4;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_A5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_A6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_AO5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_AO6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_A_CY;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_A_XOR;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_B;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_B1;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_B2;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_B3;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_B4;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_B5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_B6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_BO5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_BO6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_B_CY;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_B_XOR;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_C;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_C1;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_C2;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_C3;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_C4;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_C5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_C6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_CO5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_CO6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_C_CY;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_C_XOR;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_D;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_D1;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_D2;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_D3;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_D4;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_D5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_D6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_DO5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_DO6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_D_CY;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X14Y5_D_XOR;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_A;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_A1;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_A2;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_A3;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_A4;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_A5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_A6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_AMUX;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_AO5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_AO6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_AQ;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_AX;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_A_CY;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_A_XOR;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_B;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_B1;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_B2;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_B3;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_B4;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_B5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_B6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_BMUX;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_BO5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_BO6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_BQ;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_BX;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_B_CY;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_B_XOR;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_C;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_C1;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_C2;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_C3;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_C4;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_C5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_C6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_CLK;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_CMUX;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_CO5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_CO6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_COUT;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_CQ;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_CX;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_C_CY;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_C_XOR;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_D;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_D1;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_D2;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_D3;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_D4;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_D5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_D6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_DMUX;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_DO5;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_DO6;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_DQ;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_DX;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_D_CY;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_D_XOR;
  wire [0:0] CLBLM_R_X11Y5_SLICE_X15Y5_SR;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_A;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_A1;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_A2;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_A3;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_A4;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_A5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_A6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_AO5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_AO6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_A_CY;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_A_XOR;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_B;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_B1;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_B2;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_B3;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_B4;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_B5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_B6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_BO5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_BO6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_B_CY;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_B_XOR;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_C;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_C1;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_C2;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_C3;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_C4;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_C5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_C6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_CO5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_CO6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_C_CY;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_C_XOR;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_D;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_D1;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_D2;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_D3;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_D4;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_D5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_D6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_DO5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_DO6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_D_CY;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X14Y6_D_XOR;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_A;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_A1;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_A2;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_A3;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_A4;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_A5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_A6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_AMUX;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_AO5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_AO6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_AQ;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_AX;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_A_CY;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_A_XOR;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_B;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_B1;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_B2;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_B3;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_B4;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_B5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_B6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_BMUX;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_BO5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_BO6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_BQ;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_BX;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_B_CY;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_B_XOR;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_C;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_C1;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_C2;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_C3;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_C4;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_C5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_C6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_CIN;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_CLK;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_CMUX;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_CO5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_CO6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_COUT;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_CQ;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_CX;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_C_CY;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_C_XOR;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_D;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_D1;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_D2;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_D3;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_D4;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_D5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_D6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_DMUX;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_DO5;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_DO6;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_DQ;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_DX;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_D_CY;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_D_XOR;
  wire [0:0] CLBLM_R_X11Y6_SLICE_X15Y6_SR;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_A;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_A1;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_A2;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_A3;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_A4;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_A5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_A6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_AO5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_AO6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_A_CY;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_A_XOR;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_B;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_B1;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_B2;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_B3;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_B4;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_B5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_B6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_BO5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_BO6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_B_CY;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_B_XOR;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_C;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_C1;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_C2;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_C3;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_C4;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_C5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_C6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_CO5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_CO6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_C_CY;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_C_XOR;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_D;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_D1;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_D2;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_D3;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_D4;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_D5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_D6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_DO5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_DO6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_D_CY;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X14Y7_D_XOR;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_A;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_A1;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_A2;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_A3;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_A4;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_A5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_A6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_AMUX;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_AO5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_AO6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_AQ;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_AX;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_A_CY;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_A_XOR;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_B;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_B1;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_B2;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_B3;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_B4;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_B5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_B6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_BMUX;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_BO5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_BO6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_BQ;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_BX;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_B_CY;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_B_XOR;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_C;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_C1;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_C2;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_C3;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_C4;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_C5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_C6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_CIN;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_CLK;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_CMUX;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_CO5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_CO6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_COUT;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_CQ;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_CX;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_C_CY;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_C_XOR;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_D;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_D1;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_D2;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_D3;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_D4;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_D5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_D6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_DMUX;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_DO5;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_DO6;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_DQ;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_DX;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_D_CY;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_D_XOR;
  wire [0:0] CLBLM_R_X11Y7_SLICE_X15Y7_SR;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_A;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_A1;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_A2;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_A3;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_A4;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_A5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_A6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_AO5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_AO6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_A_CY;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_A_XOR;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_B;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_B1;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_B2;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_B3;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_B4;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_B5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_B6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_BO5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_BO6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_B_CY;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_B_XOR;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_C;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_C1;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_C2;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_C3;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_C4;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_C5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_C6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_CO5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_CO6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_C_CY;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_C_XOR;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_D;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_D1;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_D2;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_D3;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_D4;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_D5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_D6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_DO5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_DO6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_D_CY;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X14Y8_D_XOR;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_A;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_A1;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_A2;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_A3;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_A4;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_A5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_A6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_AO5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_AO6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_AQ;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_AX;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_A_CY;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_A_XOR;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_B;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_B1;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_B2;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_B3;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_B4;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_B5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_B6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_BMUX;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_BO5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_BO6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_BQ;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_BX;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_B_CY;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_B_XOR;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_C;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_C1;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_C2;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_C3;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_C4;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_C5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_C6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_CIN;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_CLK;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_CMUX;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_CO5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_CO6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_COUT;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_CQ;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_CX;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_C_CY;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_C_XOR;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_D;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_D1;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_D2;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_D3;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_D4;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_D5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_D6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_DMUX;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_DO5;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_DO6;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_DQ;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_DX;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_D_CY;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_D_XOR;
  wire [0:0] CLBLM_R_X11Y8_SLICE_X15Y8_SR;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_A;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_A1;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_A2;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_A3;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_A4;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_A5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_A6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_AO5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_AO6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_A_CY;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_A_XOR;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_B;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_B1;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_B2;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_B3;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_B4;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_B5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_B6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_BO5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_BO6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_B_CY;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_B_XOR;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_C;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_C1;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_C2;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_C3;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_C4;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_C5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_C6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_CO5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_CO6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_C_CY;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_C_XOR;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_D;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_D1;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_D2;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_D3;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_D4;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_D5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_D6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_DO5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_DO6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_D_CY;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X14Y9_D_XOR;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_A;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_A1;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_A2;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_A3;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_A4;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_A5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_A6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_AO5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_AO6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_AQ;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_AX;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_A_CY;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_A_XOR;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_B;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_B1;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_B2;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_B3;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_B4;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_B5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_B6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_BMUX;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_BO5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_BO6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_BQ;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_BX;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_B_CY;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_B_XOR;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_C;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_C1;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_C2;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_C3;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_C4;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_C5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_C6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_CIN;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_CLK;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_CMUX;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_CO5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_CO6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_COUT;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_CQ;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_CX;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_C_CY;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_C_XOR;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_D;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_D1;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_D2;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_D3;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_D4;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_D5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_D6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_DMUX;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_DO5;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_DO6;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_DQ;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_DX;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_D_CY;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_D_XOR;
  wire [0:0] CLBLM_R_X11Y9_SLICE_X15Y9_SR;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_A;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_A1;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_A2;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_A3;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_A4;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_A5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_A6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_AO5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_AO6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_A_CY;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_A_XOR;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_B;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_B1;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_B2;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_B3;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_B4;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_B5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_B6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_BO5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_BO6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_B_CY;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_B_XOR;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_C;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_C1;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_C2;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_C3;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_C4;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_C5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_C6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_CO5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_CO6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_C_CY;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_C_XOR;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_D;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_D1;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_D2;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_D3;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_D4;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_D5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_D6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_DO5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_DO6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_D_CY;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X42Y14_D_XOR;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_A;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_A1;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_A2;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_A3;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_A4;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_A5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_A6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_AMUX;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_AO5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_AO6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_AQ;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_AX;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_A_CY;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_A_XOR;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_B;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_B1;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_B2;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_B3;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_B4;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_B5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_B6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_BMUX;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_BO5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_BO6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_BQ;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_BX;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_B_CY;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_B_XOR;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_C;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_C1;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_C2;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_C3;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_C4;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_C5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_C6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_CLK;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_CMUX;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_CO5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_CO6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_COUT;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_CQ;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_CX;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_C_CY;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_C_XOR;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_D;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_D1;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_D2;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_D3;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_D4;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_D5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_D6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_DMUX;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_DO5;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_DO6;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_DQ;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_DX;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_D_CY;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_D_XOR;
  wire [0:0] CLBLM_R_X27Y14_SLICE_X43Y14_SR;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_A;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_A1;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_A2;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_A3;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_A4;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_A5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_A6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_AO5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_AO6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_A_CY;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_A_XOR;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_B;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_B1;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_B2;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_B3;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_B4;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_B5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_B6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_BO5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_BO6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_B_CY;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_B_XOR;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_C;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_C1;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_C2;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_C3;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_C4;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_C5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_C6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_CO5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_CO6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_C_CY;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_C_XOR;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_D;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_D1;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_D2;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_D3;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_D4;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_D5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_D6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_DO5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_DO6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_D_CY;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X42Y15_D_XOR;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_A;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_A1;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_A2;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_A3;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_A4;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_A5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_A6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_AMUX;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_AO5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_AO6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_AQ;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_AX;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_A_CY;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_A_XOR;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_B;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_B1;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_B2;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_B3;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_B4;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_B5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_B6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_BMUX;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_BO5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_BO6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_BQ;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_BX;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_B_CY;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_B_XOR;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_C;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_C1;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_C2;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_C3;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_C4;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_C5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_C6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_CIN;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_CLK;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_CMUX;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_CO5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_CO6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_COUT;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_CQ;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_CX;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_C_CY;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_C_XOR;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_D;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_D1;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_D2;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_D3;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_D4;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_D5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_D6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_DMUX;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_DO5;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_DO6;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_DQ;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_DX;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_D_CY;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_D_XOR;
  wire [0:0] CLBLM_R_X27Y15_SLICE_X43Y15_SR;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_A;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_A1;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_A2;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_A3;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_A4;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_A5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_A6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_AO5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_AO6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_A_CY;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_A_XOR;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_B;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_B1;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_B2;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_B3;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_B4;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_B5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_B6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_BO5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_BO6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_B_CY;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_B_XOR;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_C;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_C1;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_C2;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_C3;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_C4;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_C5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_C6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_CO5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_CO6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_C_CY;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_C_XOR;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_D;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_D1;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_D2;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_D3;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_D4;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_D5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_D6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_DO5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_DO6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_D_CY;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X42Y16_D_XOR;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_A;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_A1;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_A2;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_A3;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_A4;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_A5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_A6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_AMUX;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_AO5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_AO6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_AQ;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_AX;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_A_CY;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_A_XOR;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_B;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_B1;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_B2;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_B3;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_B4;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_B5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_B6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_BMUX;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_BO5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_BO6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_BQ;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_BX;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_B_CY;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_B_XOR;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_C;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_C1;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_C2;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_C3;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_C4;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_C5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_C6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_CIN;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_CLK;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_CMUX;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_CO5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_CO6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_COUT;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_CQ;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_CX;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_C_CY;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_C_XOR;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_D;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_D1;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_D2;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_D3;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_D4;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_D5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_D6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_DMUX;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_DO5;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_DO6;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_DQ;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_DX;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_D_CY;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_D_XOR;
  wire [0:0] CLBLM_R_X27Y16_SLICE_X43Y16_SR;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_A;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_A1;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_A2;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_A3;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_A4;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_A5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_A6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_AO5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_AO6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_A_CY;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_A_XOR;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_B;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_B1;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_B2;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_B3;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_B4;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_B5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_B6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_BO5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_BO6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_B_CY;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_B_XOR;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_C;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_C1;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_C2;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_C3;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_C4;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_C5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_C6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_CO5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_CO6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_C_CY;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_C_XOR;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_D;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_D1;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_D2;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_D3;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_D4;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_D5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_D6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_DO5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_DO6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_D_CY;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X42Y17_D_XOR;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_A;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_A1;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_A2;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_A3;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_A4;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_A5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_A6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_AO5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_AO6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_AQ;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_AX;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_A_CY;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_A_XOR;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_B;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_B1;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_B2;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_B3;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_B4;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_B5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_B6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_BMUX;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_BO5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_BO6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_BQ;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_BX;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_B_CY;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_B_XOR;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_C;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_C1;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_C2;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_C3;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_C4;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_C5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_C6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_CIN;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_CLK;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_CMUX;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_CO5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_CO6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_COUT;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_CQ;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_CX;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_C_CY;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_C_XOR;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_D;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_D1;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_D2;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_D3;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_D4;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_D5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_D6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_DMUX;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_DO5;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_DO6;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_DQ;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_DX;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_D_CY;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_D_XOR;
  wire [0:0] CLBLM_R_X27Y17_SLICE_X43Y17_SR;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_A;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_A1;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_A2;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_A3;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_A4;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_A5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_A6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_AO5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_AO6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_A_CY;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_A_XOR;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_B;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_B1;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_B2;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_B3;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_B4;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_B5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_B6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_BO5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_BO6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_B_CY;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_B_XOR;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_C;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_C1;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_C2;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_C3;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_C4;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_C5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_C6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_CO5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_CO6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_C_CY;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_C_XOR;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_D;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_D1;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_D2;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_D3;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_D4;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_D5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_D6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_DO5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_DO6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_D_CY;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X42Y18_D_XOR;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_A;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_A1;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_A2;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_A3;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_A4;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_A5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_A6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_AO5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_AO6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_AQ;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_AX;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_A_CY;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_A_XOR;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_B;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_B1;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_B2;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_B3;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_B4;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_B5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_B6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_BMUX;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_BO5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_BO6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_BQ;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_BX;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_B_CY;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_B_XOR;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_C;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_C1;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_C2;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_C3;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_C4;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_C5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_C6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_CIN;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_CLK;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_CMUX;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_CO5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_CO6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_COUT;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_CQ;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_CX;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_C_CY;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_C_XOR;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_D;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_D1;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_D2;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_D3;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_D4;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_D5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_D6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_DMUX;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_DO5;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_DO6;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_DQ;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_DX;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_D_CY;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_D_XOR;
  wire [0:0] CLBLM_R_X27Y18_SLICE_X43Y18_SR;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_A;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_A1;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_A2;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_A3;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_A4;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_A5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_A6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_AO5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_AO6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_A_CY;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_A_XOR;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_B;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_B1;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_B2;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_B3;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_B4;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_B5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_B6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_BO5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_BO6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_B_CY;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_B_XOR;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_C;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_C1;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_C2;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_C3;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_C4;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_C5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_C6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_CO5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_CO6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_C_CY;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_C_XOR;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_D;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_D1;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_D2;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_D3;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_D4;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_D5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_D6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_DO5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_DO6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_D_CY;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X42Y19_D_XOR;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_A;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_A1;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_A2;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_A3;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_A4;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_A5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_A6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_AMUX;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_AO5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_AO6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_AQ;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_AX;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_A_CY;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_A_XOR;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_B;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_B1;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_B2;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_B3;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_B4;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_B5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_B6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_BMUX;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_BO5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_BO6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_BQ;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_BX;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_B_CY;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_B_XOR;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_C;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_C1;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_C2;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_C3;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_C4;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_C5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_C6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_CIN;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_CLK;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_CMUX;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_CO6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_COUT;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_CQ;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_CX;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_C_CY;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_C_XOR;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_D;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_D1;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_D2;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_D3;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_D4;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_D5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_D6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_DO5;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_DO6;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_DQ;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_DX;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_D_CY;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_D_XOR;
  wire [0:0] CLBLM_R_X27Y19_SLICE_X43Y19_SR;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_A;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_A1;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_A2;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_A3;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_A4;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_A5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_A6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_AO5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_AO6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_A_CY;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_A_XOR;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_B;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_B1;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_B2;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_B3;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_B4;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_B5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_B6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_BO5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_BO6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_B_CY;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_B_XOR;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_C;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_C1;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_C2;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_C3;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_C4;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_C5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_C6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_CO5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_CO6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_C_CY;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_C_XOR;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_D;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_D1;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_D2;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_D3;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_D4;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_D5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_D6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_DO5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_DO6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_D_CY;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X42Y38_D_XOR;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_A;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_A1;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_A2;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_A3;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_A4;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_A5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_A6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_AMUX;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_AO5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_AO6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_AQ;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_AX;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_A_CY;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_A_XOR;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_B;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_B1;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_B2;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_B3;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_B4;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_B5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_B6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_BMUX;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_BO5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_BO6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_BQ;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_BX;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_B_CY;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_B_XOR;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_C;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_C1;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_C2;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_C3;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_C4;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_C5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_C6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_CLK;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_CMUX;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_CO5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_CO6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_COUT;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_CQ;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_CX;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_C_CY;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_C_XOR;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_D;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_D1;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_D2;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_D3;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_D4;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_D5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_D6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_DMUX;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_DO5;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_DO6;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_DQ;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_DX;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_D_CY;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_D_XOR;
  wire [0:0] CLBLM_R_X27Y38_SLICE_X43Y38_SR;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_A;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_A1;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_A2;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_A3;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_A4;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_A5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_A6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_AO5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_AO6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_A_CY;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_A_XOR;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_B;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_B1;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_B2;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_B3;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_B4;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_B5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_B6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_BO5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_BO6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_B_CY;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_B_XOR;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_C;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_C1;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_C2;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_C3;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_C4;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_C5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_C6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_CO5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_CO6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_C_CY;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_C_XOR;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_D;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_D1;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_D2;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_D3;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_D4;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_D5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_D6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_DO5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_DO6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_D_CY;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X42Y39_D_XOR;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_A;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_A1;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_A2;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_A3;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_A4;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_A5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_A6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_AMUX;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_AO5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_AO6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_AQ;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_AX;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_A_CY;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_A_XOR;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_B;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_B1;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_B2;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_B3;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_B4;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_B5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_B6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_BMUX;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_BO5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_BO6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_BQ;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_BX;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_B_CY;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_B_XOR;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_C;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_C1;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_C2;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_C3;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_C4;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_C5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_C6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_CIN;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_CLK;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_CMUX;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_CO5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_CO6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_COUT;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_CQ;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_CX;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_C_CY;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_C_XOR;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_D;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_D1;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_D2;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_D3;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_D4;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_D5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_D6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_DMUX;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_DO5;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_DO6;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_DQ;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_DX;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_D_CY;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_D_XOR;
  wire [0:0] CLBLM_R_X27Y39_SLICE_X43Y39_SR;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_A;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_A1;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_A2;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_A3;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_A4;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_A5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_A6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_AO5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_AO6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_A_CY;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_A_XOR;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_B;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_B1;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_B2;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_B3;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_B4;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_B5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_B6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_BO5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_BO6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_B_CY;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_B_XOR;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_C;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_C1;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_C2;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_C3;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_C4;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_C5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_C6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_CO5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_CO6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_C_CY;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_C_XOR;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_D;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_D1;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_D2;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_D3;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_D4;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_D5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_D6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_DO5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_DO6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_D_CY;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X42Y40_D_XOR;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_A;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_A1;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_A2;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_A3;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_A4;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_A5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_A6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_AMUX;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_AO5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_AO6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_AQ;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_AX;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_A_CY;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_A_XOR;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_B;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_B1;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_B2;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_B3;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_B4;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_B5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_B6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_BMUX;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_BO5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_BO6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_BQ;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_BX;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_B_CY;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_B_XOR;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_C;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_C1;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_C2;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_C3;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_C4;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_C5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_C6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_CIN;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_CLK;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_CMUX;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_CO5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_CO6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_COUT;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_CQ;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_CX;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_C_CY;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_C_XOR;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_D;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_D1;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_D2;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_D3;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_D4;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_D5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_D6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_DMUX;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_DO5;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_DO6;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_DQ;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_DX;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_D_CY;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_D_XOR;
  wire [0:0] CLBLM_R_X27Y40_SLICE_X43Y40_SR;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_A;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_A1;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_A2;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_A3;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_A4;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_A5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_A6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_AO5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_AO6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_A_CY;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_A_XOR;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_B;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_B1;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_B2;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_B3;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_B4;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_B5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_B6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_BO5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_BO6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_B_CY;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_B_XOR;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_C;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_C1;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_C2;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_C3;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_C4;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_C5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_C6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_CO5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_CO6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_C_CY;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_C_XOR;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_D;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_D1;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_D2;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_D3;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_D4;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_D5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_D6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_DO5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_DO6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_D_CY;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X42Y41_D_XOR;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_A;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_A1;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_A2;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_A3;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_A4;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_A5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_A5Q;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_A6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_AMUX;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_AO5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_AO6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_AQ;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_AX;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_A_CY;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_A_XOR;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_B;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_B1;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_B2;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_B3;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_B4;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_B5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_B6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_BMUX;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_BO5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_BO6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_BQ;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_BX;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_B_CY;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_B_XOR;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_C;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_C1;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_C2;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_C3;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_C4;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_C5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_C6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_CIN;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_CLK;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_CMUX;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_CO5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_CO6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_COUT;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_CQ;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_CX;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_C_CY;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_C_XOR;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_D;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_D1;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_D2;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_D3;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_D4;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_D5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_D6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_DMUX;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_DO5;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_DO6;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_DQ;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_DX;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_D_CY;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_D_XOR;
  wire [0:0] CLBLM_R_X27Y41_SLICE_X43Y41_SR;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_A;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_A1;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_A2;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_A3;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_A4;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_A5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_A6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_AO5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_AO6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_A_CY;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_A_XOR;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_B;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_B1;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_B2;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_B3;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_B4;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_B5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_B6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_BO5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_BO6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_B_CY;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_B_XOR;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_C;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_C1;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_C2;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_C3;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_C4;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_C5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_C6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_CO5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_CO6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_C_CY;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_C_XOR;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_D;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_D1;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_D2;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_D3;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_D4;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_D5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_D6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_DO5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_DO6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_D_CY;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X42Y42_D_XOR;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_A;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_A1;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_A2;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_A3;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_A4;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_A5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_A5Q;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_A6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_AMUX;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_AO5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_AO6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_AQ;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_AX;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_A_CY;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_A_XOR;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_B;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_B1;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_B2;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_B3;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_B4;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_B5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_B6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_BMUX;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_BO5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_BO6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_BQ;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_BX;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_B_CY;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_B_XOR;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_C;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_C1;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_C2;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_C3;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_C4;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_C5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_C6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_CIN;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_CLK;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_CMUX;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_CO5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_CO6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_COUT;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_CQ;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_CX;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_C_CY;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_C_XOR;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_D;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_D1;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_D2;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_D3;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_D4;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_D5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_D6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_DMUX;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_DO5;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_DO6;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_DQ;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_DX;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_D_CY;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_D_XOR;
  wire [0:0] CLBLM_R_X27Y42_SLICE_X43Y42_SR;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_A;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_A1;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_A2;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_A3;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_A4;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_A5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_A6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_AO5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_AO6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_A_CY;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_A_XOR;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_B;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_B1;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_B2;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_B3;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_B4;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_B5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_B6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_BO5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_BO6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_B_CY;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_B_XOR;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_C;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_C1;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_C2;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_C3;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_C4;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_C5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_C6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_CO5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_CO6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_C_CY;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_C_XOR;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_D;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_D1;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_D2;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_D3;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_D4;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_D5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_D6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_DO5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_DO6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_D_CY;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X42Y43_D_XOR;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_A;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_A1;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_A2;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_A3;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_A4;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_A5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_A6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_AMUX;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_AO5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_AO6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_AX;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_A_CY;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_A_XOR;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_B;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_B1;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_B2;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_B3;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_B4;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_B5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_B6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_BMUX;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_BO5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_BO6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_BX;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_B_CY;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_B_XOR;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_C;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_C1;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_C2;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_C3;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_C4;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_C5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_C6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_CIN;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_CLK;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_CMUX;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_CO5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_CO6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_COUT;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_CQ;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_CX;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_C_CY;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_C_XOR;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_D;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_D1;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_D2;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_D3;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_D4;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_D5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_D6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_DMUX;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_DO5;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_DO6;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_DQ;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_DX;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_D_CY;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_D_XOR;
  wire [0:0] CLBLM_R_X27Y43_SLICE_X43Y43_SR;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_A;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_A1;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_A2;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_A3;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_A4;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_A5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_A6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_AO5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_AO6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_A_CY;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_A_XOR;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_B;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_B1;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_B2;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_B3;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_B4;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_B5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_B6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_BO5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_BO6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_BQ;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_BX;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_B_CY;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_B_XOR;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_C;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_C1;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_C2;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_C3;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_C4;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_C5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_C6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_CLK;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_CO5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_CO6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_CQ;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_CX;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_C_CY;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_C_XOR;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_D;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_D1;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_D2;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_D3;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_D4;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_D5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_D6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_DO5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_DO6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_DQ;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_DX;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_D_CY;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_D_XOR;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X42Y8_SR;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_A;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_A1;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_A2;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_A3;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_A4;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_A5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_A6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_AO5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_AO6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_A_CY;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_A_XOR;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_B;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_B1;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_B2;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_B3;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_B4;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_B5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_B6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_BO5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_BO6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_B_CY;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_B_XOR;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_C;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_C1;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_C2;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_C3;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_C4;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_C5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_C6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_CO5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_CO6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_C_CY;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_C_XOR;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_D;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_D1;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_D2;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_D3;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_D4;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_D5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_D6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_DO5;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_DO6;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_D_CY;
  wire [0:0] CLBLM_R_X27Y8_SLICE_X43Y8_D_XOR;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_A;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_A1;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_A2;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_A3;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_A4;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_A5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_A6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_AMUX;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_AO5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_AO6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_AX;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_A_CY;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_A_XOR;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_B;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_B1;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_B2;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_B3;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_B4;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_B5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_B6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_BMUX;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_BO5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_BO6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_BX;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_B_CY;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_B_XOR;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_C;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_C1;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_C2;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_C3;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_C4;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_C5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_C6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_CIN;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_CLK;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_CMUX;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_CO5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_CO6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_COUT;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_CQ;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_CX;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_C_CY;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_C_XOR;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_D;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_D1;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_D2;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_D3;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_D4;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_D5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_D6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_DMUX;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_DO5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_DO6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_DQ;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_DX;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_D_CY;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_D_XOR;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X2Y10_SR;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_A;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_A1;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_A2;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_A3;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_A4;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_A5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_A6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_AO5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_AO6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_A_CY;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_A_XOR;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_B;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_B1;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_B2;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_B3;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_B4;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_B5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_B6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_BO5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_BO6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_B_CY;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_B_XOR;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_C;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_C1;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_C2;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_C3;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_C4;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_C5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_C6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_CO5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_CO6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_C_CY;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_C_XOR;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_D;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_D1;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_D2;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_D3;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_D4;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_D5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_D6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_DO5;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_DO6;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_D_CY;
  wire [0:0] CLBLM_R_X3Y10_SLICE_X3Y10_D_XOR;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_A;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_A1;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_A2;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_A3;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_A4;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_A5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_A6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_AMUX;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_AO5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_AO6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_AQ;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_AX;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_A_CY;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_A_XOR;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_B;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_B1;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_B2;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_B3;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_B4;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_B5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_B6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_BMUX;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_BO5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_BO6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_BQ;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_BX;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_B_CY;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_B_XOR;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_C;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_C1;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_C2;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_C3;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_C4;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_C5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_C6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_CLK;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_CMUX;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_CO5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_CO6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_COUT;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_CQ;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_CX;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_C_CY;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_C_XOR;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_D;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_D1;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_D2;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_D3;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_D4;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_D5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_D6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_DMUX;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_DO5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_DO6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_DQ;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_DX;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_D_CY;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_D_XOR;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X2Y5_SR;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_A;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_A1;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_A2;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_A3;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_A4;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_A5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_A6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_AO5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_AO6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_A_CY;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_A_XOR;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_B;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_B1;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_B2;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_B3;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_B4;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_B5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_B6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_BO5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_BO6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_B_CY;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_B_XOR;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_C;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_C1;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_C2;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_C3;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_C4;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_C5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_C6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_CO5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_CO6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_C_CY;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_C_XOR;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_D;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_D1;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_D2;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_D3;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_D4;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_D5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_D6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_DO5;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_DO6;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_D_CY;
  wire [0:0] CLBLM_R_X3Y5_SLICE_X3Y5_D_XOR;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_A;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_A1;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_A2;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_A3;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_A4;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_A5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_A6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_AMUX;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_AO5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_AO6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_AQ;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_AX;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_A_CY;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_A_XOR;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_B;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_B1;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_B2;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_B3;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_B4;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_B5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_B6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_BMUX;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_BO5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_BO6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_BQ;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_BX;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_B_CY;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_B_XOR;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_C;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_C1;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_C2;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_C3;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_C4;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_C5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_C6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_CIN;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_CLK;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_CMUX;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_CO5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_CO6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_COUT;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_CQ;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_CX;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_C_CY;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_C_XOR;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_D;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_D1;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_D2;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_D3;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_D4;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_D5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_D6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_DMUX;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_DO5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_DO6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_DQ;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_DX;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_D_CY;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_D_XOR;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X2Y6_SR;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_A;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_A1;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_A2;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_A3;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_A4;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_A5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_A6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_AO5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_AO6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_A_CY;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_A_XOR;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_B;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_B1;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_B2;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_B3;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_B4;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_B5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_B6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_BO5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_BO6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_B_CY;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_B_XOR;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_C;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_C1;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_C2;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_C3;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_C4;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_C5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_C6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_CO5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_CO6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_C_CY;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_C_XOR;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_D;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_D1;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_D2;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_D3;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_D4;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_D5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_D6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_DO5;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_DO6;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_D_CY;
  wire [0:0] CLBLM_R_X3Y6_SLICE_X3Y6_D_XOR;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_A;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_A1;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_A2;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_A3;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_A4;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_A5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_A6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_AMUX;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_AO5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_AO6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_AQ;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_AX;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_A_CY;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_A_XOR;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_B;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_B1;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_B2;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_B3;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_B4;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_B5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_B6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_BMUX;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_BO5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_BO6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_BQ;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_BX;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_B_CY;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_B_XOR;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_C;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_C1;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_C2;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_C3;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_C4;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_C5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_C6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_CIN;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_CLK;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_CMUX;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_CO5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_CO6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_COUT;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_CQ;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_CX;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_C_CY;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_C_XOR;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_D;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_D1;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_D2;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_D3;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_D4;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_D5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_D6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_DMUX;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_DO5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_DO6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_DQ;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_DX;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_D_CY;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_D_XOR;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X2Y7_SR;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_A;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_A1;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_A2;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_A3;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_A4;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_A5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_A6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_AO5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_AO6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_A_CY;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_A_XOR;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_B;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_B1;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_B2;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_B3;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_B4;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_B5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_B6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_BO5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_BO6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_B_CY;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_B_XOR;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_C;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_C1;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_C2;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_C3;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_C4;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_C5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_C6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_CO5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_CO6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_C_CY;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_C_XOR;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_D;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_D1;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_D2;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_D3;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_D4;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_D5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_D6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_DO5;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_DO6;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_D_CY;
  wire [0:0] CLBLM_R_X3Y7_SLICE_X3Y7_D_XOR;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_A;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_A1;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_A2;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_A3;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_A4;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_A5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_A5Q;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_A6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_AMUX;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_AO5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_AO6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_AQ;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_AX;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_A_CY;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_A_XOR;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_B;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_B1;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_B2;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_B3;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_B4;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_B5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_B6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_BMUX;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_BO5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_BO6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_BQ;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_BX;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_B_CY;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_B_XOR;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_C;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_C1;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_C2;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_C3;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_C4;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_C5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_C6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_CIN;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_CLK;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_CMUX;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_CO5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_CO6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_COUT;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_CQ;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_CX;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_C_CY;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_C_XOR;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_D;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_D1;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_D2;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_D3;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_D4;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_D5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_D6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_DMUX;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_DO5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_DO6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_DQ;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_DX;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_D_CY;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_D_XOR;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X2Y8_SR;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_A;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_A1;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_A2;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_A3;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_A4;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_A5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_A6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_AO5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_AO6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_A_CY;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_A_XOR;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_B;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_B1;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_B2;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_B3;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_B4;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_B5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_B6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_BO5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_BO6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_B_CY;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_B_XOR;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_C;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_C1;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_C2;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_C3;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_C4;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_C5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_C6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_CO5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_CO6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_C_CY;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_C_XOR;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_D;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_D1;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_D2;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_D3;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_D4;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_D5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_D6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_DO5;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_DO6;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_D_CY;
  wire [0:0] CLBLM_R_X3Y8_SLICE_X3Y8_D_XOR;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_A;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_A1;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_A2;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_A3;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_A4;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_A5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_A6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_AMUX;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_AO5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_AO6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_AQ;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_AX;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_A_CY;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_A_XOR;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_B;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_B1;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_B2;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_B3;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_B4;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_B5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_B6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_BMUX;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_BO5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_BO6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_BQ;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_BX;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_B_CY;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_B_XOR;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_C;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_C1;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_C2;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_C3;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_C4;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_C5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_C5Q;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_C6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_CIN;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_CLK;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_CMUX;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_CO5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_CO6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_COUT;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_CQ;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_CX;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_C_CY;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_C_XOR;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_D;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_D1;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_D2;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_D3;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_D4;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_D5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_D6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_DMUX;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_DO5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_DO6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_DQ;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_DX;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_D_CY;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_D_XOR;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X2Y9_SR;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_A;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_A1;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_A2;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_A3;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_A4;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_A5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_A6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_AO5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_AO6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_A_CY;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_A_XOR;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_B;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_B1;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_B2;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_B3;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_B4;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_B5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_B6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_BO5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_BO6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_B_CY;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_B_XOR;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_C;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_C1;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_C2;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_C3;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_C4;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_C5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_C6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_CO5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_CO6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_C_CY;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_C_XOR;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_D;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_D1;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_D2;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_D3;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_D4;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_D5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_D6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_DO5;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_DO6;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_D_CY;
  wire [0:0] CLBLM_R_X3Y9_SLICE_X3Y9_D_XOR;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_A;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_A1;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_A2;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_A3;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_A4;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_A5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_A6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_AO5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_AO6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_A_CY;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_A_XOR;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_B;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_B1;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_B2;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_B3;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_B4;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_B5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_B6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_BO5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_BO6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_B_CY;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_B_XOR;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_C;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_C1;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_C2;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_C3;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_C4;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_C5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_C6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_CO5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_CO6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_C_CY;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_C_XOR;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_D;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_D1;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_D2;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_D3;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_D4;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_D5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_D6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_DO5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_DO6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_D_CY;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X6Y15_D_XOR;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_A;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_A1;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_A2;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_A3;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_A4;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_A5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_A6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_AMUX;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_AO5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_AO6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_AQ;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_AX;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_A_CY;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_A_XOR;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_B;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_B1;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_B2;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_B3;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_B4;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_B5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_B6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_BMUX;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_BO5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_BO6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_BQ;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_BX;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_B_CY;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_B_XOR;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_C;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_C1;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_C2;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_C3;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_C4;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_C5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_C6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_CLK;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_CMUX;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_CO5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_CO6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_COUT;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_CQ;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_CX;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_C_CY;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_C_XOR;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_D;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_D1;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_D2;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_D3;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_D4;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_D5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_D6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_DMUX;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_DO5;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_DO6;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_DQ;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_DX;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_D_CY;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_D_XOR;
  wire [0:0] CLBLM_R_X5Y15_SLICE_X7Y15_SR;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_A;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_A1;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_A2;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_A3;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_A4;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_A5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_A6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_AO5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_AO6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_A_CY;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_A_XOR;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_B;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_B1;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_B2;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_B3;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_B4;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_B5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_B6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_BO5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_BO6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_B_CY;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_B_XOR;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_C;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_C1;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_C2;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_C3;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_C4;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_C5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_C6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_CO5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_CO6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_C_CY;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_C_XOR;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_D;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_D1;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_D2;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_D3;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_D4;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_D5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_D6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_DO5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_DO6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_D_CY;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X6Y16_D_XOR;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_A;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_A1;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_A2;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_A3;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_A4;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_A5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_A6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_AMUX;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_AO5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_AO6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_AQ;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_AX;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_A_CY;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_A_XOR;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_B;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_B1;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_B2;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_B3;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_B4;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_B5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_B6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_BMUX;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_BO5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_BO6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_BQ;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_BX;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_B_CY;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_B_XOR;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_C;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_C1;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_C2;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_C3;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_C4;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_C5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_C6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_CIN;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_CLK;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_CMUX;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_CO5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_CO6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_COUT;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_CQ;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_CX;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_C_CY;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_C_XOR;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_D;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_D1;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_D2;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_D3;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_D4;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_D5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_D6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_DMUX;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_DO5;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_DO6;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_DQ;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_DX;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_D_CY;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_D_XOR;
  wire [0:0] CLBLM_R_X5Y16_SLICE_X7Y16_SR;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_A;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_A1;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_A2;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_A3;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_A4;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_A5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_A6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_AO5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_AO6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_A_CY;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_A_XOR;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_B;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_B1;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_B2;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_B3;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_B4;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_B5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_B6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_BO5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_BO6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_B_CY;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_B_XOR;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_C;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_C1;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_C2;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_C3;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_C4;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_C5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_C6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_CO5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_CO6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_C_CY;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_C_XOR;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_D;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_D1;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_D2;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_D3;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_D4;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_D5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_D6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_DO5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_DO6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_D_CY;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X6Y17_D_XOR;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_A;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_A1;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_A2;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_A3;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_A4;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_A5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_A6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_AMUX;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_AO5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_AO6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_AQ;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_AX;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_A_CY;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_A_XOR;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_B;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_B1;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_B2;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_B3;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_B4;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_B5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_B6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_BMUX;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_BO5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_BO6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_BQ;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_BX;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_B_CY;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_B_XOR;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_C;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_C1;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_C2;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_C3;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_C4;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_C5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_C6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_CIN;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_CLK;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_CMUX;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_CO5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_CO6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_COUT;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_CQ;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_CX;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_C_CY;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_C_XOR;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_D;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_D1;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_D2;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_D3;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_D4;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_D5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_D6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_DMUX;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_DO5;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_DO6;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_DQ;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_DX;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_D_CY;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_D_XOR;
  wire [0:0] CLBLM_R_X5Y17_SLICE_X7Y17_SR;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_A;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_A1;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_A2;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_A3;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_A4;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_A5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_A6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_AO5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_AO6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_A_CY;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_A_XOR;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_B;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_B1;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_B2;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_B3;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_B4;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_B5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_B6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_BO5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_BO6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_B_CY;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_B_XOR;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_C;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_C1;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_C2;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_C3;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_C4;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_C5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_C6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_CO5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_CO6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_C_CY;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_C_XOR;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_D;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_D1;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_D2;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_D3;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_D4;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_D5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_D6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_DO5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_DO6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_D_CY;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X6Y18_D_XOR;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_A;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_A1;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_A2;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_A3;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_A4;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_A5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_A6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_AO5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_AO6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_AQ;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_AX;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_A_CY;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_A_XOR;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_B;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_B1;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_B2;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_B3;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_B4;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_B5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_B6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_BMUX;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_BO5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_BO6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_BQ;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_BX;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_B_CY;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_B_XOR;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_C;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_C1;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_C2;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_C3;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_C4;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_C5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_C6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_CIN;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_CLK;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_CMUX;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_CO5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_CO6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_COUT;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_CQ;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_CX;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_C_CY;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_C_XOR;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_D;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_D1;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_D2;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_D3;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_D4;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_D5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_D6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_DMUX;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_DO5;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_DO6;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_DQ;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_DX;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_D_CY;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_D_XOR;
  wire [0:0] CLBLM_R_X5Y18_SLICE_X7Y18_SR;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_A;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_A1;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_A2;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_A3;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_A4;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_A5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_A6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_AO5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_AO6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_A_CY;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_A_XOR;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_B;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_B1;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_B2;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_B3;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_B4;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_B5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_B6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_BO5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_BO6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_B_CY;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_B_XOR;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_C;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_C1;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_C2;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_C3;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_C4;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_C5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_C6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_CO5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_CO6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_C_CY;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_C_XOR;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_D;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_D1;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_D2;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_D3;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_D4;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_D5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_D6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_DO5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_DO6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_D_CY;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X6Y19_D_XOR;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_A;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_A1;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_A2;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_A3;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_A4;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_A5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_A6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_AO5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_AO6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_AQ;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_AX;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_A_CY;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_A_XOR;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_B;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_B1;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_B2;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_B3;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_B4;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_B5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_B6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_BMUX;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_BO5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_BO6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_BQ;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_BX;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_B_CY;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_B_XOR;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_C;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_C1;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_C2;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_C3;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_C4;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_C5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_C6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_CIN;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_CLK;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_CMUX;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_CO5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_CO6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_COUT;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_CQ;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_CX;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_C_CY;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_C_XOR;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_D;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_D1;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_D2;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_D3;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_D4;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_D5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_D6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_DMUX;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_DO5;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_DO6;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_DQ;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_DX;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_D_CY;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_D_XOR;
  wire [0:0] CLBLM_R_X5Y19_SLICE_X7Y19_SR;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_A;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_A1;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_A2;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_A3;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_A4;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_A5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_A6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_AO5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_AO6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_A_CY;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_A_XOR;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_B;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_B1;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_B2;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_B3;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_B4;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_B5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_B6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_BO5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_BO6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_B_CY;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_B_XOR;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_C;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_C1;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_C2;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_C3;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_C4;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_C5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_C6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_CO5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_CO6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_C_CY;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_C_XOR;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_D;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_D1;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_D2;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_D3;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_D4;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_D5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_D6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_DO5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_DO6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_D_CY;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X6Y20_D_XOR;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_A;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_A1;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_A2;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_A3;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_A4;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_A5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_A6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_AMUX;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_AO5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_AO6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_AQ;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_AX;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_A_CY;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_A_XOR;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_B;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_B1;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_B2;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_B3;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_B4;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_B5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_B6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_BMUX;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_BO5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_BO6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_BQ;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_BX;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_B_CY;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_B_XOR;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_C;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_C1;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_C2;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_C3;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_C4;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_C5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_C6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_CIN;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_CLK;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_CO5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_CO6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_COUT;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_CQ;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_CX;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_C_CY;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_C_XOR;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_D;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_D1;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_D2;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_D3;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_D4;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_D5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_D6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_DO5;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_DO6;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_DQ;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_DX;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_D_CY;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_D_XOR;
  wire [0:0] CLBLM_R_X5Y20_SLICE_X7Y20_SR;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_S1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_S1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_S1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_S1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_S1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_S1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S1;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_CE;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_I;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_CE;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_I;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_CE;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_I;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_CE;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_I;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_CE;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_I;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y11_CE;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y11_I;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y11_O;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_CE;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_I;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y8_CE;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y8_I;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y8_O;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBIN;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBOUT;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBOUTB;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBSTOPPED;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKIN1;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKIN2;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKINSEL;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKINSTOPPED;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT0;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT0B;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT1;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT1B;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT2;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT2B;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT3;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT3B;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT4;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT5;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR0;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR1;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR2;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR3;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR4;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR5;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR6;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DCLK;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DEN;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI0;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI1;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI10;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI11;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI12;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI13;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI14;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI15;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI2;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI3;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI4;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI5;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI6;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI7;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI8;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI9;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO0;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO1;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO10;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO11;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO12;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO13;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO14;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO15;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO2;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO3;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO4;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO5;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO6;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO7;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO8;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO9;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DRDY;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DWE;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_LOCKED;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSCLK;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSDONE;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSEN;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSINCDEC;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PWRDWN;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_RST;
  wire [0:0] LIOB33_SING_X0Y0_IOB_X0Y0_O;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y11_I;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y12_I;
  wire [0:0] LIOB33_X0Y17_IOB_X0Y18_O;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y19_O;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y20_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_O;
  wire [0:0] LIOB33_X0Y25_IOB_X0Y26_I;
  wire [0:0] LIOB33_X0Y27_IOB_X0Y28_O;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y3_O;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y4_O;
  wire [0:0] LIOB33_X0Y43_IOB_X0Y43_O;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y6_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y10_I;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_D1;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_OQ;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_T1;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_O;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_O;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_D1;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_OQ;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_T1;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_TQ;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y26_D;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y26_O;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_D1;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_OQ;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_T1;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_TQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_D1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_OQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_T1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_TQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_D1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_OQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_T1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_TQ;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_D;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_O;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_O;
  wire [0:0] RIOB33_X43Y25_IOB_X1Y26_I;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_D;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_O;


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X24Y46_SLICE_X36Y46_D_FDRE (
.C(RIOB33_X43Y25_IOB_X1Y26_I),
.CE(1'b1),
.D(CLBLL_L_X24Y46_SLICE_X36Y46_AO6),
.Q(CLBLL_L_X24Y46_SLICE_X36Y46_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X24Y46_SLICE_X36Y46_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X24Y46_SLICE_X36Y46_DO5),
.O6(CLBLL_L_X24Y46_SLICE_X36Y46_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X24Y46_SLICE_X36Y46_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X24Y46_SLICE_X36Y46_CO5),
.O6(CLBLL_L_X24Y46_SLICE_X36Y46_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X24Y46_SLICE_X36Y46_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X24Y46_SLICE_X36Y46_BO5),
.O6(CLBLL_L_X24Y46_SLICE_X36Y46_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333333300000000)
  ) CLBLL_L_X24Y46_SLICE_X36Y46_ALUT (
.I0(1'b1),
.I1(CLBLL_L_X24Y46_SLICE_X36Y46_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X24Y46_SLICE_X36Y46_AO5),
.O6(CLBLL_L_X24Y46_SLICE_X36Y46_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X24Y46_SLICE_X37Y46_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X24Y46_SLICE_X37Y46_DO5),
.O6(CLBLL_L_X24Y46_SLICE_X37Y46_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X24Y46_SLICE_X37Y46_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X24Y46_SLICE_X37Y46_CO5),
.O6(CLBLL_L_X24Y46_SLICE_X37Y46_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X24Y46_SLICE_X37Y46_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X24Y46_SLICE_X37Y46_BO5),
.O6(CLBLL_L_X24Y46_SLICE_X37Y46_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X24Y46_SLICE_X37Y46_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X24Y46_SLICE_X37Y46_AO5),
.O6(CLBLL_L_X24Y46_SLICE_X37Y46_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X26Y9_SLICE_X40Y9_D_FDRE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y11_O),
.CE(1'b1),
.D(LIOB33_X0Y11_IOB_X0Y11_I),
.Q(CLBLL_L_X26Y9_SLICE_X40Y9_DQ),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y9_SLICE_X40Y9_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y9_SLICE_X40Y9_DO5),
.O6(CLBLL_L_X26Y9_SLICE_X40Y9_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y9_SLICE_X40Y9_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y9_SLICE_X40Y9_CO5),
.O6(CLBLL_L_X26Y9_SLICE_X40Y9_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y9_SLICE_X40Y9_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y9_SLICE_X40Y9_BO5),
.O6(CLBLL_L_X26Y9_SLICE_X40Y9_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y9_SLICE_X40Y9_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y9_SLICE_X40Y9_AO5),
.O6(CLBLL_L_X26Y9_SLICE_X40Y9_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y9_SLICE_X41Y9_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y9_SLICE_X41Y9_DO5),
.O6(CLBLL_L_X26Y9_SLICE_X41Y9_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y9_SLICE_X41Y9_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y9_SLICE_X41Y9_CO5),
.O6(CLBLL_L_X26Y9_SLICE_X41Y9_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y9_SLICE_X41Y9_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y9_SLICE_X41Y9_BO5),
.O6(CLBLL_L_X26Y9_SLICE_X41Y9_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X26Y9_SLICE_X41Y9_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X26Y9_SLICE_X41Y9_AO5),
.O6(CLBLL_L_X26Y9_SLICE_X41Y9_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y5_SLICE_X2Y5_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y5_SLICE_X2Y5_AO5),
.Q(CLBLM_R_X3Y5_SLICE_X2Y5_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y5_SLICE_X2Y5_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y5_SLICE_X2Y5_BO5),
.Q(CLBLM_R_X3Y5_SLICE_X2Y5_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y5_SLICE_X2Y5_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y5_SLICE_X2Y5_CO5),
.Q(CLBLM_R_X3Y5_SLICE_X2Y5_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y5_SLICE_X2Y5_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y5_SLICE_X2Y5_DO5),
.Q(CLBLM_R_X3Y5_SLICE_X2Y5_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y5_SLICE_X2Y5_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X3Y5_SLICE_X2Y5_D_CY, CLBLM_R_X3Y5_SLICE_X2Y5_C_CY, CLBLM_R_X3Y5_SLICE_X2Y5_B_CY, CLBLM_R_X3Y5_SLICE_X2Y5_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({CLBLM_R_X3Y5_SLICE_X2Y5_D_XOR, CLBLM_R_X3Y5_SLICE_X2Y5_C_XOR, CLBLM_R_X3Y5_SLICE_X2Y5_B_XOR, CLBLM_R_X3Y5_SLICE_X2Y5_A_XOR}),
.S({CLBLM_R_X3Y5_SLICE_X2Y5_DO6, CLBLM_R_X3Y5_SLICE_X2Y5_CO6, CLBLM_R_X3Y5_SLICE_X2Y5_BO6, CLBLM_R_X3Y5_SLICE_X2Y5_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0f0f0f0)
  ) CLBLM_R_X3Y5_SLICE_X2Y5_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y5_SLICE_X2Y5_AO6),
.I3(1'b1),
.I4(CLBLM_R_X3Y5_SLICE_X2Y5_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y5_SLICE_X2Y5_DO5),
.O6(CLBLM_R_X3Y5_SLICE_X2Y5_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacccccccc)
  ) CLBLM_R_X3Y5_SLICE_X2Y5_CLUT (
.I0(CLBLM_R_X3Y5_SLICE_X2Y5_AQ),
.I1(CLBLM_R_X3Y5_SLICE_X2Y5_B_XOR),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y5_SLICE_X2Y5_CO5),
.O6(CLBLM_R_X3Y5_SLICE_X2Y5_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X3Y5_SLICE_X2Y5_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y5_SLICE_X2Y5_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y5_SLICE_X2Y5_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X3Y5_SLICE_X2Y5_BO5),
.O6(CLBLM_R_X3Y5_SLICE_X2Y5_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0fffff0000)
  ) CLBLM_R_X3Y5_SLICE_X2Y5_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y5_SLICE_X2Y5_DQ),
.I3(1'b1),
.I4(CLBLM_R_X3Y5_SLICE_X2Y5_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X3Y5_SLICE_X2Y5_AO5),
.O6(CLBLM_R_X3Y5_SLICE_X2Y5_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y5_SLICE_X3Y5_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y5_SLICE_X3Y5_DO5),
.O6(CLBLM_R_X3Y5_SLICE_X3Y5_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y5_SLICE_X3Y5_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y5_SLICE_X3Y5_CO5),
.O6(CLBLM_R_X3Y5_SLICE_X3Y5_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y5_SLICE_X3Y5_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y5_SLICE_X3Y5_BO5),
.O6(CLBLM_R_X3Y5_SLICE_X3Y5_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y5_SLICE_X3Y5_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y5_SLICE_X3Y5_AO5),
.O6(CLBLM_R_X3Y5_SLICE_X3Y5_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y6_SLICE_X2Y6_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y6_SLICE_X2Y6_AO5),
.Q(CLBLM_R_X3Y6_SLICE_X2Y6_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y6_SLICE_X2Y6_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y6_SLICE_X2Y6_BO5),
.Q(CLBLM_R_X3Y6_SLICE_X2Y6_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y6_SLICE_X2Y6_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y6_SLICE_X2Y6_CO5),
.Q(CLBLM_R_X3Y6_SLICE_X2Y6_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y6_SLICE_X2Y6_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y6_SLICE_X2Y6_DO5),
.Q(CLBLM_R_X3Y6_SLICE_X2Y6_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y6_SLICE_X2Y6_CARRY4 (
.CI(CLBLM_R_X3Y5_SLICE_X2Y5_COUT),
.CO({CLBLM_R_X3Y6_SLICE_X2Y6_D_CY, CLBLM_R_X3Y6_SLICE_X2Y6_C_CY, CLBLM_R_X3Y6_SLICE_X2Y6_B_CY, CLBLM_R_X3Y6_SLICE_X2Y6_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X3Y6_SLICE_X2Y6_D_XOR, CLBLM_R_X3Y6_SLICE_X2Y6_C_XOR, CLBLM_R_X3Y6_SLICE_X2Y6_B_XOR, CLBLM_R_X3Y6_SLICE_X2Y6_A_XOR}),
.S({CLBLM_R_X3Y6_SLICE_X2Y6_DO6, CLBLM_R_X3Y6_SLICE_X2Y6_CO6, CLBLM_R_X3Y6_SLICE_X2Y6_BO6, CLBLM_R_X3Y6_SLICE_X2Y6_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLM_R_X3Y6_SLICE_X2Y6_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y6_SLICE_X2Y6_B_XOR),
.I4(CLBLM_R_X3Y6_SLICE_X2Y6_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y6_SLICE_X2Y6_DO5),
.O6(CLBLM_R_X3Y6_SLICE_X2Y6_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X3Y6_SLICE_X2Y6_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y6_SLICE_X2Y6_A_XOR),
.I2(CLBLM_R_X3Y6_SLICE_X2Y6_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y6_SLICE_X2Y6_CO5),
.O6(CLBLM_R_X3Y6_SLICE_X2Y6_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X3Y6_SLICE_X2Y6_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y6_SLICE_X2Y6_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y6_SLICE_X2Y6_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X3Y6_SLICE_X2Y6_BO5),
.O6(CLBLM_R_X3Y6_SLICE_X2Y6_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X3Y6_SLICE_X2Y6_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y6_SLICE_X2Y6_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y6_SLICE_X2Y6_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X3Y6_SLICE_X2Y6_AO5),
.O6(CLBLM_R_X3Y6_SLICE_X2Y6_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y6_SLICE_X3Y6_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y6_SLICE_X3Y6_DO5),
.O6(CLBLM_R_X3Y6_SLICE_X3Y6_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y6_SLICE_X3Y6_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y6_SLICE_X3Y6_CO5),
.O6(CLBLM_R_X3Y6_SLICE_X3Y6_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y6_SLICE_X3Y6_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y6_SLICE_X3Y6_BO5),
.O6(CLBLM_R_X3Y6_SLICE_X3Y6_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y6_SLICE_X3Y6_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y6_SLICE_X3Y6_AO5),
.O6(CLBLM_R_X3Y6_SLICE_X3Y6_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y7_SLICE_X2Y7_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y7_SLICE_X2Y7_AO5),
.Q(CLBLM_R_X3Y7_SLICE_X2Y7_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y7_SLICE_X2Y7_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y7_SLICE_X2Y7_BO5),
.Q(CLBLM_R_X3Y7_SLICE_X2Y7_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y7_SLICE_X2Y7_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y7_SLICE_X2Y7_CO5),
.Q(CLBLM_R_X3Y7_SLICE_X2Y7_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y7_SLICE_X2Y7_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y7_SLICE_X2Y7_DO5),
.Q(CLBLM_R_X3Y7_SLICE_X2Y7_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y7_SLICE_X2Y7_CARRY4 (
.CI(CLBLM_R_X3Y6_SLICE_X2Y6_COUT),
.CO({CLBLM_R_X3Y7_SLICE_X2Y7_D_CY, CLBLM_R_X3Y7_SLICE_X2Y7_C_CY, CLBLM_R_X3Y7_SLICE_X2Y7_B_CY, CLBLM_R_X3Y7_SLICE_X2Y7_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X3Y7_SLICE_X2Y7_D_XOR, CLBLM_R_X3Y7_SLICE_X2Y7_C_XOR, CLBLM_R_X3Y7_SLICE_X2Y7_B_XOR, CLBLM_R_X3Y7_SLICE_X2Y7_A_XOR}),
.S({CLBLM_R_X3Y7_SLICE_X2Y7_DO6, CLBLM_R_X3Y7_SLICE_X2Y7_CO6, CLBLM_R_X3Y7_SLICE_X2Y7_BO6, CLBLM_R_X3Y7_SLICE_X2Y7_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLM_R_X3Y7_SLICE_X2Y7_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y7_SLICE_X2Y7_B_XOR),
.I4(CLBLM_R_X3Y7_SLICE_X2Y7_BQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y7_SLICE_X2Y7_DO5),
.O6(CLBLM_R_X3Y7_SLICE_X2Y7_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X3Y7_SLICE_X2Y7_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y7_SLICE_X2Y7_A_XOR),
.I2(CLBLM_R_X3Y7_SLICE_X2Y7_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y7_SLICE_X2Y7_CO5),
.O6(CLBLM_R_X3Y7_SLICE_X2Y7_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X3Y7_SLICE_X2Y7_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y7_SLICE_X2Y7_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y7_SLICE_X2Y7_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X3Y7_SLICE_X2Y7_BO5),
.O6(CLBLM_R_X3Y7_SLICE_X2Y7_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X3Y7_SLICE_X2Y7_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y7_SLICE_X2Y7_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y7_SLICE_X2Y7_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X3Y7_SLICE_X2Y7_AO5),
.O6(CLBLM_R_X3Y7_SLICE_X2Y7_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y7_SLICE_X3Y7_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y7_SLICE_X3Y7_DO5),
.O6(CLBLM_R_X3Y7_SLICE_X3Y7_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y7_SLICE_X3Y7_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y7_SLICE_X3Y7_CO5),
.O6(CLBLM_R_X3Y7_SLICE_X3Y7_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y7_SLICE_X3Y7_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y7_SLICE_X3Y7_BO5),
.O6(CLBLM_R_X3Y7_SLICE_X3Y7_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y7_SLICE_X3Y7_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y7_SLICE_X3Y7_AO5),
.O6(CLBLM_R_X3Y7_SLICE_X3Y7_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y8_SLICE_X2Y8_A5_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y8_SLICE_X2Y8_AO5),
.Q(CLBLM_R_X3Y8_SLICE_X2Y8_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y8_SLICE_X2Y8_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y8_SLICE_X2Y8_A_XOR),
.Q(CLBLM_R_X3Y8_SLICE_X2Y8_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y8_SLICE_X2Y8_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y8_SLICE_X2Y8_BO5),
.Q(CLBLM_R_X3Y8_SLICE_X2Y8_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y8_SLICE_X2Y8_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y8_SLICE_X2Y8_CO5),
.Q(CLBLM_R_X3Y8_SLICE_X2Y8_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y8_SLICE_X2Y8_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y8_SLICE_X2Y8_DO5),
.Q(CLBLM_R_X3Y8_SLICE_X2Y8_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y8_SLICE_X2Y8_CARRY4 (
.CI(CLBLM_R_X3Y7_SLICE_X2Y7_COUT),
.CO({CLBLM_R_X3Y8_SLICE_X2Y8_D_CY, CLBLM_R_X3Y8_SLICE_X2Y8_C_CY, CLBLM_R_X3Y8_SLICE_X2Y8_B_CY, CLBLM_R_X3Y8_SLICE_X2Y8_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X3Y8_SLICE_X2Y8_D_XOR, CLBLM_R_X3Y8_SLICE_X2Y8_C_XOR, CLBLM_R_X3Y8_SLICE_X2Y8_B_XOR, CLBLM_R_X3Y8_SLICE_X2Y8_A_XOR}),
.S({CLBLM_R_X3Y8_SLICE_X2Y8_DO6, CLBLM_R_X3Y8_SLICE_X2Y8_CO6, CLBLM_R_X3Y8_SLICE_X2Y8_BO6, CLBLM_R_X3Y8_SLICE_X2Y8_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X3Y8_SLICE_X2Y8_DLUT (
.I0(CLBLM_R_X3Y8_SLICE_X2Y8_B_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y8_SLICE_X2Y8_CQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y8_SLICE_X2Y8_DO5),
.O6(CLBLM_R_X3Y8_SLICE_X2Y8_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X3Y8_SLICE_X2Y8_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y8_SLICE_X2Y8_D_XOR),
.I2(CLBLM_R_X3Y8_SLICE_X2Y8_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y8_SLICE_X2Y8_CO5),
.O6(CLBLM_R_X3Y8_SLICE_X2Y8_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLM_R_X3Y8_SLICE_X2Y8_BLUT (
.I0(CLBLM_R_X3Y8_SLICE_X2Y8_C_XOR),
.I1(CLBLM_R_X3Y8_SLICE_X2Y8_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y8_SLICE_X2Y8_BO5),
.O6(CLBLM_R_X3Y8_SLICE_X2Y8_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0f0f0f0)
  ) CLBLM_R_X3Y8_SLICE_X2Y8_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y8_SLICE_X2Y8_AQ),
.I2(CLBLM_R_X3Y9_SLICE_X2Y9_D_XOR),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y8_SLICE_X2Y8_AO5),
.O6(CLBLM_R_X3Y8_SLICE_X2Y8_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y8_SLICE_X3Y8_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y8_SLICE_X3Y8_DO5),
.O6(CLBLM_R_X3Y8_SLICE_X3Y8_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y8_SLICE_X3Y8_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y8_SLICE_X3Y8_CO5),
.O6(CLBLM_R_X3Y8_SLICE_X3Y8_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y8_SLICE_X3Y8_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y8_SLICE_X3Y8_BO5),
.O6(CLBLM_R_X3Y8_SLICE_X3Y8_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y8_SLICE_X3Y8_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y8_SLICE_X3Y8_AO5),
.O6(CLBLM_R_X3Y8_SLICE_X3Y8_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C5FF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y9_SLICE_X2Y9_C5_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y9_SLICE_X2Y9_CO5),
.Q(CLBLM_R_X3Y9_SLICE_X2Y9_C5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y9_SLICE_X2Y9_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y9_SLICE_X2Y9_AO5),
.Q(CLBLM_R_X3Y9_SLICE_X2Y9_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y9_SLICE_X2Y9_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y9_SLICE_X2Y9_BO5),
.Q(CLBLM_R_X3Y9_SLICE_X2Y9_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y9_SLICE_X2Y9_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y9_SLICE_X2Y9_C_XOR),
.Q(CLBLM_R_X3Y9_SLICE_X2Y9_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y9_SLICE_X2Y9_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y9_SLICE_X2Y9_DO5),
.Q(CLBLM_R_X3Y9_SLICE_X2Y9_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y9_SLICE_X2Y9_CARRY4 (
.CI(CLBLM_R_X3Y8_SLICE_X2Y8_COUT),
.CO({CLBLM_R_X3Y9_SLICE_X2Y9_D_CY, CLBLM_R_X3Y9_SLICE_X2Y9_C_CY, CLBLM_R_X3Y9_SLICE_X2Y9_B_CY, CLBLM_R_X3Y9_SLICE_X2Y9_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X3Y9_SLICE_X2Y9_D_XOR, CLBLM_R_X3Y9_SLICE_X2Y9_C_XOR, CLBLM_R_X3Y9_SLICE_X2Y9_B_XOR, CLBLM_R_X3Y9_SLICE_X2Y9_A_XOR}),
.S({CLBLM_R_X3Y9_SLICE_X2Y9_DO6, CLBLM_R_X3Y9_SLICE_X2Y9_CO6, CLBLM_R_X3Y9_SLICE_X2Y9_BO6, CLBLM_R_X3Y9_SLICE_X2Y9_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X3Y9_SLICE_X2Y9_DLUT (
.I0(CLBLM_R_X3Y9_SLICE_X2Y9_B_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y8_SLICE_X2Y8_A5Q),
.I5(1'b1),
.O5(CLBLM_R_X3Y9_SLICE_X2Y9_DO5),
.O6(CLBLM_R_X3Y9_SLICE_X2Y9_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ff00)
  ) CLBLM_R_X3Y9_SLICE_X2Y9_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X3Y9_SLICE_X2Y9_CQ),
.I3(CLBLM_R_X3Y10_SLICE_X2Y10_C_XOR),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y9_SLICE_X2Y9_CO5),
.O6(CLBLM_R_X3Y9_SLICE_X2Y9_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X3Y9_SLICE_X2Y9_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y9_SLICE_X2Y9_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X3Y9_SLICE_X2Y9_A_XOR),
.I5(1'b1),
.O5(CLBLM_R_X3Y9_SLICE_X2Y9_BO5),
.O6(CLBLM_R_X3Y9_SLICE_X2Y9_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0f0f0f0)
  ) CLBLM_R_X3Y9_SLICE_X2Y9_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y9_SLICE_X2Y9_BQ),
.I2(CLBLM_R_X3Y10_SLICE_X2Y10_D_XOR),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y9_SLICE_X2Y9_AO5),
.O6(CLBLM_R_X3Y9_SLICE_X2Y9_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y9_SLICE_X3Y9_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y9_SLICE_X3Y9_DO5),
.O6(CLBLM_R_X3Y9_SLICE_X3Y9_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y9_SLICE_X3Y9_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y9_SLICE_X3Y9_CO5),
.O6(CLBLM_R_X3Y9_SLICE_X3Y9_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y9_SLICE_X3Y9_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y9_SLICE_X3Y9_BO5),
.O6(CLBLM_R_X3Y9_SLICE_X3Y9_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y9_SLICE_X3Y9_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y9_SLICE_X3Y9_AO5),
.O6(CLBLM_R_X3Y9_SLICE_X3Y9_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y10_SLICE_X2Y10_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y10_SLICE_X2Y10_CO5),
.Q(CLBLM_R_X3Y10_SLICE_X2Y10_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X3Y10_SLICE_X2Y10_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X3Y10_SLICE_X2Y10_DO5),
.Q(CLBLM_R_X3Y10_SLICE_X2Y10_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X3Y10_SLICE_X2Y10_CARRY4 (
.CI(CLBLM_R_X3Y9_SLICE_X2Y9_COUT),
.CO({CLBLM_R_X3Y10_SLICE_X2Y10_D_CY, CLBLM_R_X3Y10_SLICE_X2Y10_C_CY, CLBLM_R_X3Y10_SLICE_X2Y10_B_CY, CLBLM_R_X3Y10_SLICE_X2Y10_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X3Y10_SLICE_X2Y10_D_XOR, CLBLM_R_X3Y10_SLICE_X2Y10_C_XOR, CLBLM_R_X3Y10_SLICE_X2Y10_B_XOR, CLBLM_R_X3Y10_SLICE_X2Y10_A_XOR}),
.S({CLBLM_R_X3Y10_SLICE_X2Y10_DO6, CLBLM_R_X3Y10_SLICE_X2Y10_CO6, CLBLM_R_X3Y10_SLICE_X2Y10_BO6, CLBLM_R_X3Y10_SLICE_X2Y10_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLM_R_X3Y10_SLICE_X2Y10_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y10_SLICE_X2Y10_A_XOR),
.I4(CLBLM_R_X3Y9_SLICE_X2Y9_AQ),
.I5(1'b1),
.O5(CLBLM_R_X3Y10_SLICE_X2Y10_DO5),
.O6(CLBLM_R_X3Y10_SLICE_X2Y10_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00aaaaaaaa)
  ) CLBLM_R_X3Y10_SLICE_X2Y10_CLUT (
.I0(CLBLM_R_X3Y10_SLICE_X2Y10_B_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X3Y9_SLICE_X2Y9_C5Q),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y10_SLICE_X2Y10_CO5),
.O6(CLBLM_R_X3Y10_SLICE_X2Y10_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X3Y10_SLICE_X2Y10_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y10_SLICE_X2Y10_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y10_SLICE_X2Y10_BO5),
.O6(CLBLM_R_X3Y10_SLICE_X2Y10_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X3Y10_SLICE_X2Y10_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X3Y10_SLICE_X2Y10_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y10_SLICE_X2Y10_AO5),
.O6(CLBLM_R_X3Y10_SLICE_X2Y10_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y10_SLICE_X3Y10_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y10_SLICE_X3Y10_DO5),
.O6(CLBLM_R_X3Y10_SLICE_X3Y10_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y10_SLICE_X3Y10_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y10_SLICE_X3Y10_CO5),
.O6(CLBLM_R_X3Y10_SLICE_X3Y10_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y10_SLICE_X3Y10_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y10_SLICE_X3Y10_BO5),
.O6(CLBLM_R_X3Y10_SLICE_X3Y10_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X3Y10_SLICE_X3Y10_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X3Y10_SLICE_X3Y10_AO5),
.O6(CLBLM_R_X3Y10_SLICE_X3Y10_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y15_SLICE_X6Y15_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y15_SLICE_X6Y15_DO5),
.O6(CLBLM_R_X5Y15_SLICE_X6Y15_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y15_SLICE_X6Y15_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y15_SLICE_X6Y15_CO5),
.O6(CLBLM_R_X5Y15_SLICE_X6Y15_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y15_SLICE_X6Y15_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y15_SLICE_X6Y15_BO5),
.O6(CLBLM_R_X5Y15_SLICE_X6Y15_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y15_SLICE_X6Y15_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y15_SLICE_X6Y15_AO5),
.O6(CLBLM_R_X5Y15_SLICE_X6Y15_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y15_SLICE_X7Y15_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y15_SLICE_X7Y15_AO5),
.Q(CLBLM_R_X5Y15_SLICE_X7Y15_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y15_SLICE_X7Y15_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y15_SLICE_X7Y15_BO5),
.Q(CLBLM_R_X5Y15_SLICE_X7Y15_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y15_SLICE_X7Y15_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y15_SLICE_X7Y15_CO5),
.Q(CLBLM_R_X5Y15_SLICE_X7Y15_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y15_SLICE_X7Y15_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y15_SLICE_X7Y15_DO5),
.Q(CLBLM_R_X5Y15_SLICE_X7Y15_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y15_SLICE_X7Y15_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X5Y15_SLICE_X7Y15_D_CY, CLBLM_R_X5Y15_SLICE_X7Y15_C_CY, CLBLM_R_X5Y15_SLICE_X7Y15_B_CY, CLBLM_R_X5Y15_SLICE_X7Y15_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({CLBLM_R_X5Y15_SLICE_X7Y15_D_XOR, CLBLM_R_X5Y15_SLICE_X7Y15_C_XOR, CLBLM_R_X5Y15_SLICE_X7Y15_B_XOR, CLBLM_R_X5Y15_SLICE_X7Y15_A_XOR}),
.S({CLBLM_R_X5Y15_SLICE_X7Y15_DO6, CLBLM_R_X5Y15_SLICE_X7Y15_CO6, CLBLM_R_X5Y15_SLICE_X7Y15_BO6, CLBLM_R_X5Y15_SLICE_X7Y15_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0f0f0f0)
  ) CLBLM_R_X5Y15_SLICE_X7Y15_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y15_SLICE_X7Y15_AO6),
.I3(1'b1),
.I4(CLBLM_R_X5Y15_SLICE_X7Y15_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y15_SLICE_X7Y15_DO5),
.O6(CLBLM_R_X5Y15_SLICE_X7Y15_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacccccccc)
  ) CLBLM_R_X5Y15_SLICE_X7Y15_CLUT (
.I0(CLBLM_R_X5Y15_SLICE_X7Y15_AQ),
.I1(CLBLM_R_X5Y15_SLICE_X7Y15_B_XOR),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y15_SLICE_X7Y15_CO5),
.O6(CLBLM_R_X5Y15_SLICE_X7Y15_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X5Y15_SLICE_X7Y15_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y15_SLICE_X7Y15_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y15_SLICE_X7Y15_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X5Y15_SLICE_X7Y15_BO5),
.O6(CLBLM_R_X5Y15_SLICE_X7Y15_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0fffff0000)
  ) CLBLM_R_X5Y15_SLICE_X7Y15_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y15_SLICE_X7Y15_DQ),
.I3(1'b1),
.I4(CLBLM_R_X5Y15_SLICE_X7Y15_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X5Y15_SLICE_X7Y15_AO5),
.O6(CLBLM_R_X5Y15_SLICE_X7Y15_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y16_SLICE_X6Y16_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y16_SLICE_X6Y16_DO5),
.O6(CLBLM_R_X5Y16_SLICE_X6Y16_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y16_SLICE_X6Y16_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y16_SLICE_X6Y16_CO5),
.O6(CLBLM_R_X5Y16_SLICE_X6Y16_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y16_SLICE_X6Y16_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y16_SLICE_X6Y16_BO5),
.O6(CLBLM_R_X5Y16_SLICE_X6Y16_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y16_SLICE_X6Y16_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y16_SLICE_X6Y16_AO5),
.O6(CLBLM_R_X5Y16_SLICE_X6Y16_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y16_SLICE_X7Y16_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y16_SLICE_X7Y16_AO5),
.Q(CLBLM_R_X5Y16_SLICE_X7Y16_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y16_SLICE_X7Y16_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y16_SLICE_X7Y16_BO5),
.Q(CLBLM_R_X5Y16_SLICE_X7Y16_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y16_SLICE_X7Y16_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y16_SLICE_X7Y16_CO5),
.Q(CLBLM_R_X5Y16_SLICE_X7Y16_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y16_SLICE_X7Y16_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y16_SLICE_X7Y16_DO5),
.Q(CLBLM_R_X5Y16_SLICE_X7Y16_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y16_SLICE_X7Y16_CARRY4 (
.CI(CLBLM_R_X5Y15_SLICE_X7Y15_COUT),
.CO({CLBLM_R_X5Y16_SLICE_X7Y16_D_CY, CLBLM_R_X5Y16_SLICE_X7Y16_C_CY, CLBLM_R_X5Y16_SLICE_X7Y16_B_CY, CLBLM_R_X5Y16_SLICE_X7Y16_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X5Y16_SLICE_X7Y16_D_XOR, CLBLM_R_X5Y16_SLICE_X7Y16_C_XOR, CLBLM_R_X5Y16_SLICE_X7Y16_B_XOR, CLBLM_R_X5Y16_SLICE_X7Y16_A_XOR}),
.S({CLBLM_R_X5Y16_SLICE_X7Y16_DO6, CLBLM_R_X5Y16_SLICE_X7Y16_CO6, CLBLM_R_X5Y16_SLICE_X7Y16_BO6, CLBLM_R_X5Y16_SLICE_X7Y16_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLM_R_X5Y16_SLICE_X7Y16_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y16_SLICE_X7Y16_B_XOR),
.I4(CLBLM_R_X5Y16_SLICE_X7Y16_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y16_SLICE_X7Y16_DO5),
.O6(CLBLM_R_X5Y16_SLICE_X7Y16_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X5Y16_SLICE_X7Y16_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y16_SLICE_X7Y16_A_XOR),
.I2(CLBLM_R_X5Y16_SLICE_X7Y16_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y16_SLICE_X7Y16_CO5),
.O6(CLBLM_R_X5Y16_SLICE_X7Y16_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X5Y16_SLICE_X7Y16_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y16_SLICE_X7Y16_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y16_SLICE_X7Y16_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X5Y16_SLICE_X7Y16_BO5),
.O6(CLBLM_R_X5Y16_SLICE_X7Y16_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X5Y16_SLICE_X7Y16_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y16_SLICE_X7Y16_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y16_SLICE_X7Y16_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X5Y16_SLICE_X7Y16_AO5),
.O6(CLBLM_R_X5Y16_SLICE_X7Y16_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y17_SLICE_X6Y17_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y17_SLICE_X6Y17_DO5),
.O6(CLBLM_R_X5Y17_SLICE_X6Y17_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y17_SLICE_X6Y17_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y17_SLICE_X6Y17_CO5),
.O6(CLBLM_R_X5Y17_SLICE_X6Y17_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y17_SLICE_X6Y17_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y17_SLICE_X6Y17_BO5),
.O6(CLBLM_R_X5Y17_SLICE_X6Y17_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y17_SLICE_X6Y17_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y17_SLICE_X6Y17_AO5),
.O6(CLBLM_R_X5Y17_SLICE_X6Y17_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y17_SLICE_X7Y17_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y17_SLICE_X7Y17_AO5),
.Q(CLBLM_R_X5Y17_SLICE_X7Y17_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y17_SLICE_X7Y17_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y17_SLICE_X7Y17_BO5),
.Q(CLBLM_R_X5Y17_SLICE_X7Y17_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y17_SLICE_X7Y17_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y17_SLICE_X7Y17_CO5),
.Q(CLBLM_R_X5Y17_SLICE_X7Y17_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y17_SLICE_X7Y17_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y17_SLICE_X7Y17_DO5),
.Q(CLBLM_R_X5Y17_SLICE_X7Y17_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y17_SLICE_X7Y17_CARRY4 (
.CI(CLBLM_R_X5Y16_SLICE_X7Y16_COUT),
.CO({CLBLM_R_X5Y17_SLICE_X7Y17_D_CY, CLBLM_R_X5Y17_SLICE_X7Y17_C_CY, CLBLM_R_X5Y17_SLICE_X7Y17_B_CY, CLBLM_R_X5Y17_SLICE_X7Y17_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X5Y17_SLICE_X7Y17_D_XOR, CLBLM_R_X5Y17_SLICE_X7Y17_C_XOR, CLBLM_R_X5Y17_SLICE_X7Y17_B_XOR, CLBLM_R_X5Y17_SLICE_X7Y17_A_XOR}),
.S({CLBLM_R_X5Y17_SLICE_X7Y17_DO6, CLBLM_R_X5Y17_SLICE_X7Y17_CO6, CLBLM_R_X5Y17_SLICE_X7Y17_BO6, CLBLM_R_X5Y17_SLICE_X7Y17_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLM_R_X5Y17_SLICE_X7Y17_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X5Y17_SLICE_X7Y17_B_XOR),
.I4(CLBLM_R_X5Y17_SLICE_X7Y17_BQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y17_SLICE_X7Y17_DO5),
.O6(CLBLM_R_X5Y17_SLICE_X7Y17_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X5Y17_SLICE_X7Y17_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y17_SLICE_X7Y17_A_XOR),
.I2(CLBLM_R_X5Y17_SLICE_X7Y17_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y17_SLICE_X7Y17_CO5),
.O6(CLBLM_R_X5Y17_SLICE_X7Y17_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X5Y17_SLICE_X7Y17_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y17_SLICE_X7Y17_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y17_SLICE_X7Y17_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X5Y17_SLICE_X7Y17_BO5),
.O6(CLBLM_R_X5Y17_SLICE_X7Y17_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X5Y17_SLICE_X7Y17_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y17_SLICE_X7Y17_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y17_SLICE_X7Y17_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X5Y17_SLICE_X7Y17_AO5),
.O6(CLBLM_R_X5Y17_SLICE_X7Y17_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y18_SLICE_X6Y18_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y18_SLICE_X6Y18_DO5),
.O6(CLBLM_R_X5Y18_SLICE_X6Y18_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y18_SLICE_X6Y18_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y18_SLICE_X6Y18_CO5),
.O6(CLBLM_R_X5Y18_SLICE_X6Y18_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y18_SLICE_X6Y18_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y18_SLICE_X6Y18_BO5),
.O6(CLBLM_R_X5Y18_SLICE_X6Y18_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y18_SLICE_X6Y18_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y18_SLICE_X6Y18_AO5),
.O6(CLBLM_R_X5Y18_SLICE_X6Y18_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y18_SLICE_X7Y18_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y18_SLICE_X7Y18_A_XOR),
.Q(CLBLM_R_X5Y18_SLICE_X7Y18_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y18_SLICE_X7Y18_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y18_SLICE_X7Y18_BO5),
.Q(CLBLM_R_X5Y18_SLICE_X7Y18_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y18_SLICE_X7Y18_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y18_SLICE_X7Y18_CO5),
.Q(CLBLM_R_X5Y18_SLICE_X7Y18_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y18_SLICE_X7Y18_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y18_SLICE_X7Y18_DO5),
.Q(CLBLM_R_X5Y18_SLICE_X7Y18_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y18_SLICE_X7Y18_CARRY4 (
.CI(CLBLM_R_X5Y17_SLICE_X7Y17_COUT),
.CO({CLBLM_R_X5Y18_SLICE_X7Y18_D_CY, CLBLM_R_X5Y18_SLICE_X7Y18_C_CY, CLBLM_R_X5Y18_SLICE_X7Y18_B_CY, CLBLM_R_X5Y18_SLICE_X7Y18_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X5Y18_SLICE_X7Y18_D_XOR, CLBLM_R_X5Y18_SLICE_X7Y18_C_XOR, CLBLM_R_X5Y18_SLICE_X7Y18_B_XOR, CLBLM_R_X5Y18_SLICE_X7Y18_A_XOR}),
.S({CLBLM_R_X5Y18_SLICE_X7Y18_DO6, CLBLM_R_X5Y18_SLICE_X7Y18_CO6, CLBLM_R_X5Y18_SLICE_X7Y18_BO6, CLBLM_R_X5Y18_SLICE_X7Y18_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X5Y18_SLICE_X7Y18_DLUT (
.I0(CLBLM_R_X5Y18_SLICE_X7Y18_B_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y18_SLICE_X7Y18_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y18_SLICE_X7Y18_DO5),
.O6(CLBLM_R_X5Y18_SLICE_X7Y18_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X5Y18_SLICE_X7Y18_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y18_SLICE_X7Y18_D_XOR),
.I2(CLBLM_R_X5Y18_SLICE_X7Y18_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y18_SLICE_X7Y18_CO5),
.O6(CLBLM_R_X5Y18_SLICE_X7Y18_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLM_R_X5Y18_SLICE_X7Y18_BLUT (
.I0(CLBLM_R_X5Y18_SLICE_X7Y18_C_XOR),
.I1(CLBLM_R_X5Y18_SLICE_X7Y18_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y18_SLICE_X7Y18_BO5),
.O6(CLBLM_R_X5Y18_SLICE_X7Y18_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X5Y18_SLICE_X7Y18_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y18_SLICE_X7Y18_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y18_SLICE_X7Y18_AO5),
.O6(CLBLM_R_X5Y18_SLICE_X7Y18_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y19_SLICE_X6Y19_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y19_SLICE_X6Y19_DO5),
.O6(CLBLM_R_X5Y19_SLICE_X6Y19_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y19_SLICE_X6Y19_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y19_SLICE_X6Y19_CO5),
.O6(CLBLM_R_X5Y19_SLICE_X6Y19_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y19_SLICE_X6Y19_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y19_SLICE_X6Y19_BO5),
.O6(CLBLM_R_X5Y19_SLICE_X6Y19_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y19_SLICE_X6Y19_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y19_SLICE_X6Y19_AO5),
.O6(CLBLM_R_X5Y19_SLICE_X6Y19_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y19_SLICE_X7Y19_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y19_SLICE_X7Y19_A_XOR),
.Q(CLBLM_R_X5Y19_SLICE_X7Y19_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y19_SLICE_X7Y19_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y19_SLICE_X7Y19_BO5),
.Q(CLBLM_R_X5Y19_SLICE_X7Y19_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y19_SLICE_X7Y19_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y19_SLICE_X7Y19_CO5),
.Q(CLBLM_R_X5Y19_SLICE_X7Y19_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y19_SLICE_X7Y19_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y19_SLICE_X7Y19_DO5),
.Q(CLBLM_R_X5Y19_SLICE_X7Y19_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y19_SLICE_X7Y19_CARRY4 (
.CI(CLBLM_R_X5Y18_SLICE_X7Y18_COUT),
.CO({CLBLM_R_X5Y19_SLICE_X7Y19_D_CY, CLBLM_R_X5Y19_SLICE_X7Y19_C_CY, CLBLM_R_X5Y19_SLICE_X7Y19_B_CY, CLBLM_R_X5Y19_SLICE_X7Y19_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X5Y19_SLICE_X7Y19_D_XOR, CLBLM_R_X5Y19_SLICE_X7Y19_C_XOR, CLBLM_R_X5Y19_SLICE_X7Y19_B_XOR, CLBLM_R_X5Y19_SLICE_X7Y19_A_XOR}),
.S({CLBLM_R_X5Y19_SLICE_X7Y19_DO6, CLBLM_R_X5Y19_SLICE_X7Y19_CO6, CLBLM_R_X5Y19_SLICE_X7Y19_BO6, CLBLM_R_X5Y19_SLICE_X7Y19_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X5Y19_SLICE_X7Y19_DLUT (
.I0(CLBLM_R_X5Y19_SLICE_X7Y19_B_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y19_SLICE_X7Y19_CQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y19_SLICE_X7Y19_DO5),
.O6(CLBLM_R_X5Y19_SLICE_X7Y19_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X5Y19_SLICE_X7Y19_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y19_SLICE_X7Y19_D_XOR),
.I2(CLBLM_R_X5Y19_SLICE_X7Y19_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y19_SLICE_X7Y19_CO5),
.O6(CLBLM_R_X5Y19_SLICE_X7Y19_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLM_R_X5Y19_SLICE_X7Y19_BLUT (
.I0(CLBLM_R_X5Y19_SLICE_X7Y19_C_XOR),
.I1(CLBLM_R_X5Y19_SLICE_X7Y19_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y19_SLICE_X7Y19_BO5),
.O6(CLBLM_R_X5Y19_SLICE_X7Y19_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X5Y19_SLICE_X7Y19_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y19_SLICE_X7Y19_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y19_SLICE_X7Y19_AO5),
.O6(CLBLM_R_X5Y19_SLICE_X7Y19_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y20_SLICE_X6Y20_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y20_SLICE_X6Y20_DO5),
.O6(CLBLM_R_X5Y20_SLICE_X6Y20_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y20_SLICE_X6Y20_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y20_SLICE_X6Y20_CO5),
.O6(CLBLM_R_X5Y20_SLICE_X6Y20_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y20_SLICE_X6Y20_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y20_SLICE_X6Y20_BO5),
.O6(CLBLM_R_X5Y20_SLICE_X6Y20_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X5Y20_SLICE_X6Y20_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y20_SLICE_X6Y20_AO5),
.O6(CLBLM_R_X5Y20_SLICE_X6Y20_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y20_SLICE_X7Y20_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y20_SLICE_X7Y20_AO5),
.Q(CLBLM_R_X5Y20_SLICE_X7Y20_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y20_SLICE_X7Y20_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y20_SLICE_X7Y20_BO5),
.Q(CLBLM_R_X5Y20_SLICE_X7Y20_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y20_SLICE_X7Y20_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y20_SLICE_X7Y20_C_XOR),
.Q(CLBLM_R_X5Y20_SLICE_X7Y20_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X5Y20_SLICE_X7Y20_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X5Y20_SLICE_X7Y20_D_XOR),
.Q(CLBLM_R_X5Y20_SLICE_X7Y20_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X5Y20_SLICE_X7Y20_CARRY4 (
.CI(CLBLM_R_X5Y19_SLICE_X7Y19_COUT),
.CO({CLBLM_R_X5Y20_SLICE_X7Y20_D_CY, CLBLM_R_X5Y20_SLICE_X7Y20_C_CY, CLBLM_R_X5Y20_SLICE_X7Y20_B_CY, CLBLM_R_X5Y20_SLICE_X7Y20_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X5Y20_SLICE_X7Y20_D_XOR, CLBLM_R_X5Y20_SLICE_X7Y20_C_XOR, CLBLM_R_X5Y20_SLICE_X7Y20_B_XOR, CLBLM_R_X5Y20_SLICE_X7Y20_A_XOR}),
.S({CLBLM_R_X5Y20_SLICE_X7Y20_DO6, CLBLM_R_X5Y20_SLICE_X7Y20_CO6, CLBLM_R_X5Y20_SLICE_X7Y20_BO6, CLBLM_R_X5Y20_SLICE_X7Y20_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000000000)
  ) CLBLM_R_X5Y20_SLICE_X7Y20_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y20_SLICE_X7Y20_DQ),
.I5(1'b1),
.O5(CLBLM_R_X5Y20_SLICE_X7Y20_DO5),
.O6(CLBLM_R_X5Y20_SLICE_X7Y20_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLM_R_X5Y20_SLICE_X7Y20_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X5Y20_SLICE_X7Y20_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X5Y20_SLICE_X7Y20_CO5),
.O6(CLBLM_R_X5Y20_SLICE_X7Y20_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X5Y20_SLICE_X7Y20_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y20_SLICE_X7Y20_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y20_SLICE_X7Y20_A_XOR),
.I5(1'b1),
.O5(CLBLM_R_X5Y20_SLICE_X7Y20_BO5),
.O6(CLBLM_R_X5Y20_SLICE_X7Y20_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X5Y20_SLICE_X7Y20_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X5Y20_SLICE_X7Y20_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X5Y20_SLICE_X7Y20_B_XOR),
.I5(1'b1),
.O5(CLBLM_R_X5Y20_SLICE_X7Y20_AO5),
.O6(CLBLM_R_X5Y20_SLICE_X7Y20_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y5_SLICE_X14Y5_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y5_SLICE_X14Y5_DO5),
.O6(CLBLM_R_X11Y5_SLICE_X14Y5_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y5_SLICE_X14Y5_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y5_SLICE_X14Y5_CO5),
.O6(CLBLM_R_X11Y5_SLICE_X14Y5_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y5_SLICE_X14Y5_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y5_SLICE_X14Y5_BO5),
.O6(CLBLM_R_X11Y5_SLICE_X14Y5_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y5_SLICE_X14Y5_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y5_SLICE_X14Y5_AO5),
.O6(CLBLM_R_X11Y5_SLICE_X14Y5_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y5_SLICE_X15Y5_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y5_SLICE_X15Y5_AO5),
.Q(CLBLM_R_X11Y5_SLICE_X15Y5_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y5_SLICE_X15Y5_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y5_SLICE_X15Y5_BO5),
.Q(CLBLM_R_X11Y5_SLICE_X15Y5_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y5_SLICE_X15Y5_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y5_SLICE_X15Y5_CO5),
.Q(CLBLM_R_X11Y5_SLICE_X15Y5_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y5_SLICE_X15Y5_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y5_SLICE_X15Y5_DO5),
.Q(CLBLM_R_X11Y5_SLICE_X15Y5_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y5_SLICE_X15Y5_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X11Y5_SLICE_X15Y5_D_CY, CLBLM_R_X11Y5_SLICE_X15Y5_C_CY, CLBLM_R_X11Y5_SLICE_X15Y5_B_CY, CLBLM_R_X11Y5_SLICE_X15Y5_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({CLBLM_R_X11Y5_SLICE_X15Y5_D_XOR, CLBLM_R_X11Y5_SLICE_X15Y5_C_XOR, CLBLM_R_X11Y5_SLICE_X15Y5_B_XOR, CLBLM_R_X11Y5_SLICE_X15Y5_A_XOR}),
.S({CLBLM_R_X11Y5_SLICE_X15Y5_DO6, CLBLM_R_X11Y5_SLICE_X15Y5_CO6, CLBLM_R_X11Y5_SLICE_X15Y5_BO6, CLBLM_R_X11Y5_SLICE_X15Y5_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0f0f0f0)
  ) CLBLM_R_X11Y5_SLICE_X15Y5_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y5_SLICE_X15Y5_AO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y5_SLICE_X15Y5_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y5_SLICE_X15Y5_DO5),
.O6(CLBLM_R_X11Y5_SLICE_X15Y5_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacccccccc)
  ) CLBLM_R_X11Y5_SLICE_X15Y5_CLUT (
.I0(CLBLM_R_X11Y5_SLICE_X15Y5_AQ),
.I1(CLBLM_R_X11Y5_SLICE_X15Y5_B_XOR),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y5_SLICE_X15Y5_CO5),
.O6(CLBLM_R_X11Y5_SLICE_X15Y5_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X11Y5_SLICE_X15Y5_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y5_SLICE_X15Y5_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y5_SLICE_X15Y5_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y5_SLICE_X15Y5_BO5),
.O6(CLBLM_R_X11Y5_SLICE_X15Y5_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0fffff0000)
  ) CLBLM_R_X11Y5_SLICE_X15Y5_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y5_SLICE_X15Y5_DQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y5_SLICE_X15Y5_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y5_SLICE_X15Y5_AO5),
.O6(CLBLM_R_X11Y5_SLICE_X15Y5_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y6_SLICE_X14Y6_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y6_SLICE_X14Y6_DO5),
.O6(CLBLM_R_X11Y6_SLICE_X14Y6_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y6_SLICE_X14Y6_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y6_SLICE_X14Y6_CO5),
.O6(CLBLM_R_X11Y6_SLICE_X14Y6_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y6_SLICE_X14Y6_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y6_SLICE_X14Y6_BO5),
.O6(CLBLM_R_X11Y6_SLICE_X14Y6_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y6_SLICE_X14Y6_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y6_SLICE_X14Y6_AO5),
.O6(CLBLM_R_X11Y6_SLICE_X14Y6_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y6_SLICE_X15Y6_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y6_SLICE_X15Y6_AO5),
.Q(CLBLM_R_X11Y6_SLICE_X15Y6_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y6_SLICE_X15Y6_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y6_SLICE_X15Y6_BO5),
.Q(CLBLM_R_X11Y6_SLICE_X15Y6_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y6_SLICE_X15Y6_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y6_SLICE_X15Y6_CO5),
.Q(CLBLM_R_X11Y6_SLICE_X15Y6_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y6_SLICE_X15Y6_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y6_SLICE_X15Y6_DO5),
.Q(CLBLM_R_X11Y6_SLICE_X15Y6_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y6_SLICE_X15Y6_CARRY4 (
.CI(CLBLM_R_X11Y5_SLICE_X15Y5_COUT),
.CO({CLBLM_R_X11Y6_SLICE_X15Y6_D_CY, CLBLM_R_X11Y6_SLICE_X15Y6_C_CY, CLBLM_R_X11Y6_SLICE_X15Y6_B_CY, CLBLM_R_X11Y6_SLICE_X15Y6_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y6_SLICE_X15Y6_D_XOR, CLBLM_R_X11Y6_SLICE_X15Y6_C_XOR, CLBLM_R_X11Y6_SLICE_X15Y6_B_XOR, CLBLM_R_X11Y6_SLICE_X15Y6_A_XOR}),
.S({CLBLM_R_X11Y6_SLICE_X15Y6_DO6, CLBLM_R_X11Y6_SLICE_X15Y6_CO6, CLBLM_R_X11Y6_SLICE_X15Y6_BO6, CLBLM_R_X11Y6_SLICE_X15Y6_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLM_R_X11Y6_SLICE_X15Y6_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y6_SLICE_X15Y6_B_XOR),
.I4(CLBLM_R_X11Y6_SLICE_X15Y6_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y6_SLICE_X15Y6_DO5),
.O6(CLBLM_R_X11Y6_SLICE_X15Y6_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X11Y6_SLICE_X15Y6_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y6_SLICE_X15Y6_A_XOR),
.I2(CLBLM_R_X11Y6_SLICE_X15Y6_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y6_SLICE_X15Y6_CO5),
.O6(CLBLM_R_X11Y6_SLICE_X15Y6_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X11Y6_SLICE_X15Y6_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y6_SLICE_X15Y6_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y6_SLICE_X15Y6_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y6_SLICE_X15Y6_BO5),
.O6(CLBLM_R_X11Y6_SLICE_X15Y6_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X11Y6_SLICE_X15Y6_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y6_SLICE_X15Y6_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y6_SLICE_X15Y6_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y6_SLICE_X15Y6_AO5),
.O6(CLBLM_R_X11Y6_SLICE_X15Y6_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y7_SLICE_X14Y7_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y7_SLICE_X14Y7_DO5),
.O6(CLBLM_R_X11Y7_SLICE_X14Y7_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y7_SLICE_X14Y7_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y7_SLICE_X14Y7_CO5),
.O6(CLBLM_R_X11Y7_SLICE_X14Y7_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y7_SLICE_X14Y7_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y7_SLICE_X14Y7_BO5),
.O6(CLBLM_R_X11Y7_SLICE_X14Y7_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y7_SLICE_X14Y7_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y7_SLICE_X14Y7_AO5),
.O6(CLBLM_R_X11Y7_SLICE_X14Y7_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y7_SLICE_X15Y7_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y7_SLICE_X15Y7_AO5),
.Q(CLBLM_R_X11Y7_SLICE_X15Y7_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y7_SLICE_X15Y7_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y7_SLICE_X15Y7_BO5),
.Q(CLBLM_R_X11Y7_SLICE_X15Y7_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y7_SLICE_X15Y7_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y7_SLICE_X15Y7_CO5),
.Q(CLBLM_R_X11Y7_SLICE_X15Y7_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y7_SLICE_X15Y7_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y7_SLICE_X15Y7_DO5),
.Q(CLBLM_R_X11Y7_SLICE_X15Y7_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y7_SLICE_X15Y7_CARRY4 (
.CI(CLBLM_R_X11Y6_SLICE_X15Y6_COUT),
.CO({CLBLM_R_X11Y7_SLICE_X15Y7_D_CY, CLBLM_R_X11Y7_SLICE_X15Y7_C_CY, CLBLM_R_X11Y7_SLICE_X15Y7_B_CY, CLBLM_R_X11Y7_SLICE_X15Y7_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y7_SLICE_X15Y7_D_XOR, CLBLM_R_X11Y7_SLICE_X15Y7_C_XOR, CLBLM_R_X11Y7_SLICE_X15Y7_B_XOR, CLBLM_R_X11Y7_SLICE_X15Y7_A_XOR}),
.S({CLBLM_R_X11Y7_SLICE_X15Y7_DO6, CLBLM_R_X11Y7_SLICE_X15Y7_CO6, CLBLM_R_X11Y7_SLICE_X15Y7_BO6, CLBLM_R_X11Y7_SLICE_X15Y7_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLM_R_X11Y7_SLICE_X15Y7_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y7_SLICE_X15Y7_B_XOR),
.I4(CLBLM_R_X11Y7_SLICE_X15Y7_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y7_SLICE_X15Y7_DO5),
.O6(CLBLM_R_X11Y7_SLICE_X15Y7_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X11Y7_SLICE_X15Y7_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y7_SLICE_X15Y7_A_XOR),
.I2(CLBLM_R_X11Y7_SLICE_X15Y7_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y7_SLICE_X15Y7_CO5),
.O6(CLBLM_R_X11Y7_SLICE_X15Y7_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X11Y7_SLICE_X15Y7_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y7_SLICE_X15Y7_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y7_SLICE_X15Y7_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y7_SLICE_X15Y7_BO5),
.O6(CLBLM_R_X11Y7_SLICE_X15Y7_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X11Y7_SLICE_X15Y7_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y7_SLICE_X15Y7_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y7_SLICE_X15Y7_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y7_SLICE_X15Y7_AO5),
.O6(CLBLM_R_X11Y7_SLICE_X15Y7_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y8_SLICE_X14Y8_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y8_SLICE_X14Y8_DO5),
.O6(CLBLM_R_X11Y8_SLICE_X14Y8_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y8_SLICE_X14Y8_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y8_SLICE_X14Y8_CO5),
.O6(CLBLM_R_X11Y8_SLICE_X14Y8_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y8_SLICE_X14Y8_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y8_SLICE_X14Y8_BO5),
.O6(CLBLM_R_X11Y8_SLICE_X14Y8_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y8_SLICE_X14Y8_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y8_SLICE_X14Y8_AO5),
.O6(CLBLM_R_X11Y8_SLICE_X14Y8_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y8_SLICE_X15Y8_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y8_SLICE_X15Y8_A_XOR),
.Q(CLBLM_R_X11Y8_SLICE_X15Y8_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y8_SLICE_X15Y8_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y8_SLICE_X15Y8_BO5),
.Q(CLBLM_R_X11Y8_SLICE_X15Y8_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y8_SLICE_X15Y8_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y8_SLICE_X15Y8_CO5),
.Q(CLBLM_R_X11Y8_SLICE_X15Y8_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y8_SLICE_X15Y8_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y8_SLICE_X15Y8_DO5),
.Q(CLBLM_R_X11Y8_SLICE_X15Y8_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y8_SLICE_X15Y8_CARRY4 (
.CI(CLBLM_R_X11Y7_SLICE_X15Y7_COUT),
.CO({CLBLM_R_X11Y8_SLICE_X15Y8_D_CY, CLBLM_R_X11Y8_SLICE_X15Y8_C_CY, CLBLM_R_X11Y8_SLICE_X15Y8_B_CY, CLBLM_R_X11Y8_SLICE_X15Y8_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y8_SLICE_X15Y8_D_XOR, CLBLM_R_X11Y8_SLICE_X15Y8_C_XOR, CLBLM_R_X11Y8_SLICE_X15Y8_B_XOR, CLBLM_R_X11Y8_SLICE_X15Y8_A_XOR}),
.S({CLBLM_R_X11Y8_SLICE_X15Y8_DO6, CLBLM_R_X11Y8_SLICE_X15Y8_CO6, CLBLM_R_X11Y8_SLICE_X15Y8_BO6, CLBLM_R_X11Y8_SLICE_X15Y8_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X11Y8_SLICE_X15Y8_DLUT (
.I0(CLBLM_R_X11Y8_SLICE_X15Y8_B_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y8_SLICE_X15Y8_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y8_SLICE_X15Y8_DO5),
.O6(CLBLM_R_X11Y8_SLICE_X15Y8_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X11Y8_SLICE_X15Y8_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y8_SLICE_X15Y8_D_XOR),
.I2(CLBLM_R_X11Y8_SLICE_X15Y8_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y8_SLICE_X15Y8_CO5),
.O6(CLBLM_R_X11Y8_SLICE_X15Y8_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLM_R_X11Y8_SLICE_X15Y8_BLUT (
.I0(CLBLM_R_X11Y8_SLICE_X15Y8_C_XOR),
.I1(CLBLM_R_X11Y8_SLICE_X15Y8_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y8_SLICE_X15Y8_BO5),
.O6(CLBLM_R_X11Y8_SLICE_X15Y8_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X11Y8_SLICE_X15Y8_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y8_SLICE_X15Y8_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y8_SLICE_X15Y8_AO5),
.O6(CLBLM_R_X11Y8_SLICE_X15Y8_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y9_SLICE_X14Y9_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y9_SLICE_X14Y9_DO5),
.O6(CLBLM_R_X11Y9_SLICE_X14Y9_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y9_SLICE_X14Y9_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y9_SLICE_X14Y9_CO5),
.O6(CLBLM_R_X11Y9_SLICE_X14Y9_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y9_SLICE_X14Y9_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y9_SLICE_X14Y9_BO5),
.O6(CLBLM_R_X11Y9_SLICE_X14Y9_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y9_SLICE_X14Y9_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y9_SLICE_X14Y9_AO5),
.O6(CLBLM_R_X11Y9_SLICE_X14Y9_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y9_SLICE_X15Y9_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y9_SLICE_X15Y9_A_XOR),
.Q(CLBLM_R_X11Y9_SLICE_X15Y9_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y9_SLICE_X15Y9_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y9_SLICE_X15Y9_BO5),
.Q(CLBLM_R_X11Y9_SLICE_X15Y9_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y9_SLICE_X15Y9_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y9_SLICE_X15Y9_CO5),
.Q(CLBLM_R_X11Y9_SLICE_X15Y9_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y9_SLICE_X15Y9_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y9_SLICE_X15Y9_DO5),
.Q(CLBLM_R_X11Y9_SLICE_X15Y9_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y9_SLICE_X15Y9_CARRY4 (
.CI(CLBLM_R_X11Y8_SLICE_X15Y8_COUT),
.CO({CLBLM_R_X11Y9_SLICE_X15Y9_D_CY, CLBLM_R_X11Y9_SLICE_X15Y9_C_CY, CLBLM_R_X11Y9_SLICE_X15Y9_B_CY, CLBLM_R_X11Y9_SLICE_X15Y9_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y9_SLICE_X15Y9_D_XOR, CLBLM_R_X11Y9_SLICE_X15Y9_C_XOR, CLBLM_R_X11Y9_SLICE_X15Y9_B_XOR, CLBLM_R_X11Y9_SLICE_X15Y9_A_XOR}),
.S({CLBLM_R_X11Y9_SLICE_X15Y9_DO6, CLBLM_R_X11Y9_SLICE_X15Y9_CO6, CLBLM_R_X11Y9_SLICE_X15Y9_BO6, CLBLM_R_X11Y9_SLICE_X15Y9_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X11Y9_SLICE_X15Y9_DLUT (
.I0(CLBLM_R_X11Y9_SLICE_X15Y9_B_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y9_SLICE_X15Y9_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y9_SLICE_X15Y9_DO5),
.O6(CLBLM_R_X11Y9_SLICE_X15Y9_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X11Y9_SLICE_X15Y9_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y9_SLICE_X15Y9_D_XOR),
.I2(CLBLM_R_X11Y9_SLICE_X15Y9_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y9_SLICE_X15Y9_CO5),
.O6(CLBLM_R_X11Y9_SLICE_X15Y9_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLM_R_X11Y9_SLICE_X15Y9_BLUT (
.I0(CLBLM_R_X11Y9_SLICE_X15Y9_C_XOR),
.I1(CLBLM_R_X11Y9_SLICE_X15Y9_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y9_SLICE_X15Y9_BO5),
.O6(CLBLM_R_X11Y9_SLICE_X15Y9_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X11Y9_SLICE_X15Y9_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y9_SLICE_X15Y9_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y9_SLICE_X15Y9_AO5),
.O6(CLBLM_R_X11Y9_SLICE_X15Y9_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y10_SLICE_X14Y10_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y10_SLICE_X14Y10_DO5),
.O6(CLBLM_R_X11Y10_SLICE_X14Y10_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y10_SLICE_X14Y10_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y10_SLICE_X14Y10_CO5),
.O6(CLBLM_R_X11Y10_SLICE_X14Y10_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y10_SLICE_X14Y10_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y10_SLICE_X14Y10_BO5),
.O6(CLBLM_R_X11Y10_SLICE_X14Y10_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y10_SLICE_X14Y10_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y10_SLICE_X14Y10_AO5),
.O6(CLBLM_R_X11Y10_SLICE_X14Y10_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y10_SLICE_X15Y10_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y10_SLICE_X15Y10_AO5),
.Q(CLBLM_R_X11Y10_SLICE_X15Y10_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y10_SLICE_X15Y10_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y10_SLICE_X15Y10_BO5),
.Q(CLBLM_R_X11Y10_SLICE_X15Y10_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y10_SLICE_X15Y10_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y10_SLICE_X15Y10_C_XOR),
.Q(CLBLM_R_X11Y10_SLICE_X15Y10_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y10_SLICE_X15Y10_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y10_SLICE_X15Y10_D_XOR),
.Q(CLBLM_R_X11Y10_SLICE_X15Y10_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y10_SLICE_X15Y10_CARRY4 (
.CI(CLBLM_R_X11Y9_SLICE_X15Y9_COUT),
.CO({CLBLM_R_X11Y10_SLICE_X15Y10_D_CY, CLBLM_R_X11Y10_SLICE_X15Y10_C_CY, CLBLM_R_X11Y10_SLICE_X15Y10_B_CY, CLBLM_R_X11Y10_SLICE_X15Y10_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y10_SLICE_X15Y10_D_XOR, CLBLM_R_X11Y10_SLICE_X15Y10_C_XOR, CLBLM_R_X11Y10_SLICE_X15Y10_B_XOR, CLBLM_R_X11Y10_SLICE_X15Y10_A_XOR}),
.S({CLBLM_R_X11Y10_SLICE_X15Y10_DO6, CLBLM_R_X11Y10_SLICE_X15Y10_CO6, CLBLM_R_X11Y10_SLICE_X15Y10_BO6, CLBLM_R_X11Y10_SLICE_X15Y10_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000000000)
  ) CLBLM_R_X11Y10_SLICE_X15Y10_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y10_SLICE_X15Y10_DQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y10_SLICE_X15Y10_DO5),
.O6(CLBLM_R_X11Y10_SLICE_X15Y10_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLM_R_X11Y10_SLICE_X15Y10_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y10_SLICE_X15Y10_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y10_SLICE_X15Y10_CO5),
.O6(CLBLM_R_X11Y10_SLICE_X15Y10_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X11Y10_SLICE_X15Y10_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y10_SLICE_X15Y10_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y10_SLICE_X15Y10_A_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y10_SLICE_X15Y10_BO5),
.O6(CLBLM_R_X11Y10_SLICE_X15Y10_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X11Y10_SLICE_X15Y10_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y10_SLICE_X15Y10_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y10_SLICE_X15Y10_B_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y10_SLICE_X15Y10_AO5),
.O6(CLBLM_R_X11Y10_SLICE_X15Y10_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y28_SLICE_X14Y28_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y28_SLICE_X14Y28_AO5),
.Q(CLBLM_R_X11Y28_SLICE_X14Y28_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y28_SLICE_X14Y28_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y28_SLICE_X14Y28_BO5),
.Q(CLBLM_R_X11Y28_SLICE_X14Y28_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y28_SLICE_X14Y28_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y28_SLICE_X14Y28_CO5),
.Q(CLBLM_R_X11Y28_SLICE_X14Y28_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y28_SLICE_X14Y28_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y28_SLICE_X14Y28_DO5),
.Q(CLBLM_R_X11Y28_SLICE_X14Y28_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y28_SLICE_X14Y28_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X11Y28_SLICE_X14Y28_D_CY, CLBLM_R_X11Y28_SLICE_X14Y28_C_CY, CLBLM_R_X11Y28_SLICE_X14Y28_B_CY, CLBLM_R_X11Y28_SLICE_X14Y28_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({CLBLM_R_X11Y28_SLICE_X14Y28_D_XOR, CLBLM_R_X11Y28_SLICE_X14Y28_C_XOR, CLBLM_R_X11Y28_SLICE_X14Y28_B_XOR, CLBLM_R_X11Y28_SLICE_X14Y28_A_XOR}),
.S({CLBLM_R_X11Y28_SLICE_X14Y28_DO6, CLBLM_R_X11Y28_SLICE_X14Y28_CO6, CLBLM_R_X11Y28_SLICE_X14Y28_BO6, CLBLM_R_X11Y28_SLICE_X14Y28_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0f0f0f0)
  ) CLBLM_R_X11Y28_SLICE_X14Y28_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y28_SLICE_X14Y28_AO6),
.I3(1'b1),
.I4(CLBLM_R_X11Y28_SLICE_X14Y28_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y28_SLICE_X14Y28_DO5),
.O6(CLBLM_R_X11Y28_SLICE_X14Y28_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacccccccc)
  ) CLBLM_R_X11Y28_SLICE_X14Y28_CLUT (
.I0(CLBLM_R_X11Y28_SLICE_X14Y28_AQ),
.I1(CLBLM_R_X11Y28_SLICE_X14Y28_B_XOR),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y28_SLICE_X14Y28_CO5),
.O6(CLBLM_R_X11Y28_SLICE_X14Y28_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X11Y28_SLICE_X14Y28_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y28_SLICE_X14Y28_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y28_SLICE_X14Y28_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y28_SLICE_X14Y28_BO5),
.O6(CLBLM_R_X11Y28_SLICE_X14Y28_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0fffff0000)
  ) CLBLM_R_X11Y28_SLICE_X14Y28_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y28_SLICE_X14Y28_DQ),
.I3(1'b1),
.I4(CLBLM_R_X11Y28_SLICE_X14Y28_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y28_SLICE_X14Y28_AO5),
.O6(CLBLM_R_X11Y28_SLICE_X14Y28_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y28_SLICE_X15Y28_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y28_SLICE_X15Y28_DO5),
.O6(CLBLM_R_X11Y28_SLICE_X15Y28_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y28_SLICE_X15Y28_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y28_SLICE_X15Y28_CO5),
.O6(CLBLM_R_X11Y28_SLICE_X15Y28_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y28_SLICE_X15Y28_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y28_SLICE_X15Y28_BO5),
.O6(CLBLM_R_X11Y28_SLICE_X15Y28_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y28_SLICE_X15Y28_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y28_SLICE_X15Y28_AO5),
.O6(CLBLM_R_X11Y28_SLICE_X15Y28_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y29_SLICE_X14Y29_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y29_SLICE_X14Y29_AO5),
.Q(CLBLM_R_X11Y29_SLICE_X14Y29_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y29_SLICE_X14Y29_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y29_SLICE_X14Y29_BO5),
.Q(CLBLM_R_X11Y29_SLICE_X14Y29_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y29_SLICE_X14Y29_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y29_SLICE_X14Y29_CO5),
.Q(CLBLM_R_X11Y29_SLICE_X14Y29_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y29_SLICE_X14Y29_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y29_SLICE_X14Y29_DO5),
.Q(CLBLM_R_X11Y29_SLICE_X14Y29_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y29_SLICE_X14Y29_CARRY4 (
.CI(CLBLM_R_X11Y28_SLICE_X14Y28_COUT),
.CO({CLBLM_R_X11Y29_SLICE_X14Y29_D_CY, CLBLM_R_X11Y29_SLICE_X14Y29_C_CY, CLBLM_R_X11Y29_SLICE_X14Y29_B_CY, CLBLM_R_X11Y29_SLICE_X14Y29_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y29_SLICE_X14Y29_D_XOR, CLBLM_R_X11Y29_SLICE_X14Y29_C_XOR, CLBLM_R_X11Y29_SLICE_X14Y29_B_XOR, CLBLM_R_X11Y29_SLICE_X14Y29_A_XOR}),
.S({CLBLM_R_X11Y29_SLICE_X14Y29_DO6, CLBLM_R_X11Y29_SLICE_X14Y29_CO6, CLBLM_R_X11Y29_SLICE_X14Y29_BO6, CLBLM_R_X11Y29_SLICE_X14Y29_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLM_R_X11Y29_SLICE_X14Y29_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y29_SLICE_X14Y29_B_XOR),
.I4(CLBLM_R_X11Y29_SLICE_X14Y29_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y29_SLICE_X14Y29_DO5),
.O6(CLBLM_R_X11Y29_SLICE_X14Y29_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X11Y29_SLICE_X14Y29_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y29_SLICE_X14Y29_A_XOR),
.I2(CLBLM_R_X11Y29_SLICE_X14Y29_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y29_SLICE_X14Y29_CO5),
.O6(CLBLM_R_X11Y29_SLICE_X14Y29_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X11Y29_SLICE_X14Y29_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y29_SLICE_X14Y29_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y29_SLICE_X14Y29_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y29_SLICE_X14Y29_BO5),
.O6(CLBLM_R_X11Y29_SLICE_X14Y29_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X11Y29_SLICE_X14Y29_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y29_SLICE_X14Y29_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y29_SLICE_X14Y29_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y29_SLICE_X14Y29_AO5),
.O6(CLBLM_R_X11Y29_SLICE_X14Y29_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y29_SLICE_X15Y29_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y29_SLICE_X15Y29_DO5),
.O6(CLBLM_R_X11Y29_SLICE_X15Y29_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y29_SLICE_X15Y29_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y29_SLICE_X15Y29_CO5),
.O6(CLBLM_R_X11Y29_SLICE_X15Y29_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y29_SLICE_X15Y29_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y29_SLICE_X15Y29_BO5),
.O6(CLBLM_R_X11Y29_SLICE_X15Y29_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y29_SLICE_X15Y29_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y29_SLICE_X15Y29_AO5),
.O6(CLBLM_R_X11Y29_SLICE_X15Y29_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y30_SLICE_X14Y30_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y30_SLICE_X14Y30_AO5),
.Q(CLBLM_R_X11Y30_SLICE_X14Y30_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y30_SLICE_X14Y30_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y30_SLICE_X14Y30_BO5),
.Q(CLBLM_R_X11Y30_SLICE_X14Y30_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y30_SLICE_X14Y30_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y30_SLICE_X14Y30_CO5),
.Q(CLBLM_R_X11Y30_SLICE_X14Y30_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y30_SLICE_X14Y30_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y30_SLICE_X14Y30_DO5),
.Q(CLBLM_R_X11Y30_SLICE_X14Y30_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y30_SLICE_X14Y30_CARRY4 (
.CI(CLBLM_R_X11Y29_SLICE_X14Y29_COUT),
.CO({CLBLM_R_X11Y30_SLICE_X14Y30_D_CY, CLBLM_R_X11Y30_SLICE_X14Y30_C_CY, CLBLM_R_X11Y30_SLICE_X14Y30_B_CY, CLBLM_R_X11Y30_SLICE_X14Y30_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y30_SLICE_X14Y30_D_XOR, CLBLM_R_X11Y30_SLICE_X14Y30_C_XOR, CLBLM_R_X11Y30_SLICE_X14Y30_B_XOR, CLBLM_R_X11Y30_SLICE_X14Y30_A_XOR}),
.S({CLBLM_R_X11Y30_SLICE_X14Y30_DO6, CLBLM_R_X11Y30_SLICE_X14Y30_CO6, CLBLM_R_X11Y30_SLICE_X14Y30_BO6, CLBLM_R_X11Y30_SLICE_X14Y30_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLM_R_X11Y30_SLICE_X14Y30_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X11Y30_SLICE_X14Y30_B_XOR),
.I4(CLBLM_R_X11Y30_SLICE_X14Y30_BQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y30_SLICE_X14Y30_DO5),
.O6(CLBLM_R_X11Y30_SLICE_X14Y30_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X11Y30_SLICE_X14Y30_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y30_SLICE_X14Y30_A_XOR),
.I2(CLBLM_R_X11Y30_SLICE_X14Y30_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y30_SLICE_X14Y30_CO5),
.O6(CLBLM_R_X11Y30_SLICE_X14Y30_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X11Y30_SLICE_X14Y30_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y30_SLICE_X14Y30_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y30_SLICE_X14Y30_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y30_SLICE_X14Y30_BO5),
.O6(CLBLM_R_X11Y30_SLICE_X14Y30_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X11Y30_SLICE_X14Y30_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y30_SLICE_X14Y30_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y30_SLICE_X14Y30_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y30_SLICE_X14Y30_AO5),
.O6(CLBLM_R_X11Y30_SLICE_X14Y30_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y30_SLICE_X15Y30_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y30_SLICE_X15Y30_DO5),
.O6(CLBLM_R_X11Y30_SLICE_X15Y30_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y30_SLICE_X15Y30_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y30_SLICE_X15Y30_CO5),
.O6(CLBLM_R_X11Y30_SLICE_X15Y30_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y30_SLICE_X15Y30_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y30_SLICE_X15Y30_BO5),
.O6(CLBLM_R_X11Y30_SLICE_X15Y30_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y30_SLICE_X15Y30_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y30_SLICE_X15Y30_AO5),
.O6(CLBLM_R_X11Y30_SLICE_X15Y30_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y31_SLICE_X14Y31_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y31_SLICE_X14Y31_A_XOR),
.Q(CLBLM_R_X11Y31_SLICE_X14Y31_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y31_SLICE_X14Y31_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y31_SLICE_X14Y31_BO5),
.Q(CLBLM_R_X11Y31_SLICE_X14Y31_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y31_SLICE_X14Y31_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y31_SLICE_X14Y31_CO5),
.Q(CLBLM_R_X11Y31_SLICE_X14Y31_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y31_SLICE_X14Y31_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y31_SLICE_X14Y31_DO5),
.Q(CLBLM_R_X11Y31_SLICE_X14Y31_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y31_SLICE_X14Y31_CARRY4 (
.CI(CLBLM_R_X11Y30_SLICE_X14Y30_COUT),
.CO({CLBLM_R_X11Y31_SLICE_X14Y31_D_CY, CLBLM_R_X11Y31_SLICE_X14Y31_C_CY, CLBLM_R_X11Y31_SLICE_X14Y31_B_CY, CLBLM_R_X11Y31_SLICE_X14Y31_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y31_SLICE_X14Y31_D_XOR, CLBLM_R_X11Y31_SLICE_X14Y31_C_XOR, CLBLM_R_X11Y31_SLICE_X14Y31_B_XOR, CLBLM_R_X11Y31_SLICE_X14Y31_A_XOR}),
.S({CLBLM_R_X11Y31_SLICE_X14Y31_DO6, CLBLM_R_X11Y31_SLICE_X14Y31_CO6, CLBLM_R_X11Y31_SLICE_X14Y31_BO6, CLBLM_R_X11Y31_SLICE_X14Y31_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X11Y31_SLICE_X14Y31_DLUT (
.I0(CLBLM_R_X11Y31_SLICE_X14Y31_B_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y31_SLICE_X14Y31_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y31_SLICE_X14Y31_DO5),
.O6(CLBLM_R_X11Y31_SLICE_X14Y31_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X11Y31_SLICE_X14Y31_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y31_SLICE_X14Y31_D_XOR),
.I2(CLBLM_R_X11Y31_SLICE_X14Y31_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y31_SLICE_X14Y31_CO5),
.O6(CLBLM_R_X11Y31_SLICE_X14Y31_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLM_R_X11Y31_SLICE_X14Y31_BLUT (
.I0(CLBLM_R_X11Y31_SLICE_X14Y31_C_XOR),
.I1(CLBLM_R_X11Y31_SLICE_X14Y31_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y31_SLICE_X14Y31_BO5),
.O6(CLBLM_R_X11Y31_SLICE_X14Y31_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X11Y31_SLICE_X14Y31_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y31_SLICE_X14Y31_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y31_SLICE_X14Y31_AO5),
.O6(CLBLM_R_X11Y31_SLICE_X14Y31_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y31_SLICE_X15Y31_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y31_SLICE_X15Y31_DO5),
.O6(CLBLM_R_X11Y31_SLICE_X15Y31_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y31_SLICE_X15Y31_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y31_SLICE_X15Y31_CO5),
.O6(CLBLM_R_X11Y31_SLICE_X15Y31_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y31_SLICE_X15Y31_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y31_SLICE_X15Y31_BO5),
.O6(CLBLM_R_X11Y31_SLICE_X15Y31_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y31_SLICE_X15Y31_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y31_SLICE_X15Y31_AO5),
.O6(CLBLM_R_X11Y31_SLICE_X15Y31_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y32_SLICE_X14Y32_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y32_SLICE_X14Y32_A_XOR),
.Q(CLBLM_R_X11Y32_SLICE_X14Y32_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y32_SLICE_X14Y32_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y32_SLICE_X14Y32_BO5),
.Q(CLBLM_R_X11Y32_SLICE_X14Y32_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y32_SLICE_X14Y32_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y32_SLICE_X14Y32_CO5),
.Q(CLBLM_R_X11Y32_SLICE_X14Y32_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y32_SLICE_X14Y32_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y32_SLICE_X14Y32_DO5),
.Q(CLBLM_R_X11Y32_SLICE_X14Y32_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y32_SLICE_X14Y32_CARRY4 (
.CI(CLBLM_R_X11Y31_SLICE_X14Y31_COUT),
.CO({CLBLM_R_X11Y32_SLICE_X14Y32_D_CY, CLBLM_R_X11Y32_SLICE_X14Y32_C_CY, CLBLM_R_X11Y32_SLICE_X14Y32_B_CY, CLBLM_R_X11Y32_SLICE_X14Y32_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y32_SLICE_X14Y32_D_XOR, CLBLM_R_X11Y32_SLICE_X14Y32_C_XOR, CLBLM_R_X11Y32_SLICE_X14Y32_B_XOR, CLBLM_R_X11Y32_SLICE_X14Y32_A_XOR}),
.S({CLBLM_R_X11Y32_SLICE_X14Y32_DO6, CLBLM_R_X11Y32_SLICE_X14Y32_CO6, CLBLM_R_X11Y32_SLICE_X14Y32_BO6, CLBLM_R_X11Y32_SLICE_X14Y32_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X11Y32_SLICE_X14Y32_DLUT (
.I0(CLBLM_R_X11Y32_SLICE_X14Y32_B_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y32_SLICE_X14Y32_CQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y32_SLICE_X14Y32_DO5),
.O6(CLBLM_R_X11Y32_SLICE_X14Y32_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X11Y32_SLICE_X14Y32_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y32_SLICE_X14Y32_D_XOR),
.I2(CLBLM_R_X11Y32_SLICE_X14Y32_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y32_SLICE_X14Y32_CO5),
.O6(CLBLM_R_X11Y32_SLICE_X14Y32_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLM_R_X11Y32_SLICE_X14Y32_BLUT (
.I0(CLBLM_R_X11Y32_SLICE_X14Y32_C_XOR),
.I1(CLBLM_R_X11Y32_SLICE_X14Y32_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y32_SLICE_X14Y32_BO5),
.O6(CLBLM_R_X11Y32_SLICE_X14Y32_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X11Y32_SLICE_X14Y32_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y32_SLICE_X14Y32_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y32_SLICE_X14Y32_AO5),
.O6(CLBLM_R_X11Y32_SLICE_X14Y32_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y32_SLICE_X15Y32_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y32_SLICE_X15Y32_DO5),
.O6(CLBLM_R_X11Y32_SLICE_X15Y32_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y32_SLICE_X15Y32_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y32_SLICE_X15Y32_CO5),
.O6(CLBLM_R_X11Y32_SLICE_X15Y32_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y32_SLICE_X15Y32_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y32_SLICE_X15Y32_BO5),
.O6(CLBLM_R_X11Y32_SLICE_X15Y32_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y32_SLICE_X15Y32_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y32_SLICE_X15Y32_AO5),
.O6(CLBLM_R_X11Y32_SLICE_X15Y32_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y33_SLICE_X14Y33_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y33_SLICE_X14Y33_AO5),
.Q(CLBLM_R_X11Y33_SLICE_X14Y33_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y33_SLICE_X14Y33_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y33_SLICE_X14Y33_BO5),
.Q(CLBLM_R_X11Y33_SLICE_X14Y33_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y33_SLICE_X14Y33_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y33_SLICE_X14Y33_C_XOR),
.Q(CLBLM_R_X11Y33_SLICE_X14Y33_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X11Y33_SLICE_X14Y33_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X11Y33_SLICE_X14Y33_D_XOR),
.Q(CLBLM_R_X11Y33_SLICE_X14Y33_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X11Y33_SLICE_X14Y33_CARRY4 (
.CI(CLBLM_R_X11Y32_SLICE_X14Y32_COUT),
.CO({CLBLM_R_X11Y33_SLICE_X14Y33_D_CY, CLBLM_R_X11Y33_SLICE_X14Y33_C_CY, CLBLM_R_X11Y33_SLICE_X14Y33_B_CY, CLBLM_R_X11Y33_SLICE_X14Y33_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X11Y33_SLICE_X14Y33_D_XOR, CLBLM_R_X11Y33_SLICE_X14Y33_C_XOR, CLBLM_R_X11Y33_SLICE_X14Y33_B_XOR, CLBLM_R_X11Y33_SLICE_X14Y33_A_XOR}),
.S({CLBLM_R_X11Y33_SLICE_X14Y33_DO6, CLBLM_R_X11Y33_SLICE_X14Y33_CO6, CLBLM_R_X11Y33_SLICE_X14Y33_BO6, CLBLM_R_X11Y33_SLICE_X14Y33_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000000000)
  ) CLBLM_R_X11Y33_SLICE_X14Y33_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y33_SLICE_X14Y33_DQ),
.I5(1'b1),
.O5(CLBLM_R_X11Y33_SLICE_X14Y33_DO5),
.O6(CLBLM_R_X11Y33_SLICE_X14Y33_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f000000000)
  ) CLBLM_R_X11Y33_SLICE_X14Y33_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X11Y33_SLICE_X14Y33_CQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y33_SLICE_X14Y33_CO5),
.O6(CLBLM_R_X11Y33_SLICE_X14Y33_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X11Y33_SLICE_X14Y33_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y33_SLICE_X14Y33_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y33_SLICE_X14Y33_A_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y33_SLICE_X14Y33_BO5),
.O6(CLBLM_R_X11Y33_SLICE_X14Y33_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X11Y33_SLICE_X14Y33_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X11Y33_SLICE_X14Y33_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X11Y33_SLICE_X14Y33_B_XOR),
.I5(1'b1),
.O5(CLBLM_R_X11Y33_SLICE_X14Y33_AO5),
.O6(CLBLM_R_X11Y33_SLICE_X14Y33_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y33_SLICE_X15Y33_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y33_SLICE_X15Y33_DO5),
.O6(CLBLM_R_X11Y33_SLICE_X15Y33_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y33_SLICE_X15Y33_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y33_SLICE_X15Y33_CO5),
.O6(CLBLM_R_X11Y33_SLICE_X15Y33_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y33_SLICE_X15Y33_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y33_SLICE_X15Y33_BO5),
.O6(CLBLM_R_X11Y33_SLICE_X15Y33_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X11Y33_SLICE_X15Y33_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X11Y33_SLICE_X15Y33_AO5),
.O6(CLBLM_R_X11Y33_SLICE_X15Y33_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y8_SLICE_X42Y8_B_FDSE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y11_O),
.CE(1'b1),
.D(CLBLL_L_X26Y9_SLICE_X40Y9_DQ),
.Q(CLBLM_R_X27Y8_SLICE_X42Y8_BQ),
.S(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y8_SLICE_X42Y8_C_FDSE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y11_O),
.CE(1'b1),
.D(CLBLM_R_X27Y8_SLICE_X42Y8_BQ),
.Q(CLBLM_R_X27Y8_SLICE_X42Y8_CQ),
.S(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDSE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y8_SLICE_X42Y8_D_FDSE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y11_O),
.CE(1'b1),
.D(CLBLM_R_X27Y8_SLICE_X42Y8_CQ),
.Q(CLBLM_R_X27Y8_SLICE_X42Y8_DQ),
.S(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y8_SLICE_X42Y8_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y8_SLICE_X42Y8_DO5),
.O6(CLBLM_R_X27Y8_SLICE_X42Y8_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y8_SLICE_X42Y8_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y8_SLICE_X42Y8_CO5),
.O6(CLBLM_R_X27Y8_SLICE_X42Y8_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y8_SLICE_X42Y8_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y8_SLICE_X42Y8_BO5),
.O6(CLBLM_R_X27Y8_SLICE_X42Y8_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y8_SLICE_X42Y8_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y8_SLICE_X42Y8_AO5),
.O6(CLBLM_R_X27Y8_SLICE_X42Y8_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y8_SLICE_X43Y8_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y8_SLICE_X43Y8_DO5),
.O6(CLBLM_R_X27Y8_SLICE_X43Y8_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y8_SLICE_X43Y8_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y8_SLICE_X43Y8_CO5),
.O6(CLBLM_R_X27Y8_SLICE_X43Y8_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y8_SLICE_X43Y8_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y8_SLICE_X43Y8_BO5),
.O6(CLBLM_R_X27Y8_SLICE_X43Y8_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y8_SLICE_X43Y8_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y8_SLICE_X43Y8_AO5),
.O6(CLBLM_R_X27Y8_SLICE_X43Y8_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y14_SLICE_X42Y14_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y14_SLICE_X42Y14_DO5),
.O6(CLBLM_R_X27Y14_SLICE_X42Y14_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y14_SLICE_X42Y14_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y14_SLICE_X42Y14_CO5),
.O6(CLBLM_R_X27Y14_SLICE_X42Y14_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y14_SLICE_X42Y14_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y14_SLICE_X42Y14_BO5),
.O6(CLBLM_R_X27Y14_SLICE_X42Y14_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y14_SLICE_X42Y14_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y14_SLICE_X42Y14_AO5),
.O6(CLBLM_R_X27Y14_SLICE_X42Y14_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y14_SLICE_X43Y14_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y14_SLICE_X43Y14_AO5),
.Q(CLBLM_R_X27Y14_SLICE_X43Y14_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y14_SLICE_X43Y14_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y14_SLICE_X43Y14_BO5),
.Q(CLBLM_R_X27Y14_SLICE_X43Y14_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y14_SLICE_X43Y14_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y14_SLICE_X43Y14_CO5),
.Q(CLBLM_R_X27Y14_SLICE_X43Y14_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y14_SLICE_X43Y14_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y14_SLICE_X43Y14_DO5),
.Q(CLBLM_R_X27Y14_SLICE_X43Y14_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X27Y14_SLICE_X43Y14_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X27Y14_SLICE_X43Y14_D_CY, CLBLM_R_X27Y14_SLICE_X43Y14_C_CY, CLBLM_R_X27Y14_SLICE_X43Y14_B_CY, CLBLM_R_X27Y14_SLICE_X43Y14_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({CLBLM_R_X27Y14_SLICE_X43Y14_D_XOR, CLBLM_R_X27Y14_SLICE_X43Y14_C_XOR, CLBLM_R_X27Y14_SLICE_X43Y14_B_XOR, CLBLM_R_X27Y14_SLICE_X43Y14_A_XOR}),
.S({CLBLM_R_X27Y14_SLICE_X43Y14_DO6, CLBLM_R_X27Y14_SLICE_X43Y14_CO6, CLBLM_R_X27Y14_SLICE_X43Y14_BO6, CLBLM_R_X27Y14_SLICE_X43Y14_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000f0f0f0f0)
  ) CLBLM_R_X27Y14_SLICE_X43Y14_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X27Y14_SLICE_X43Y14_AO6),
.I3(1'b1),
.I4(CLBLM_R_X27Y14_SLICE_X43Y14_BQ),
.I5(1'b1),
.O5(CLBLM_R_X27Y14_SLICE_X43Y14_DO5),
.O6(CLBLM_R_X27Y14_SLICE_X43Y14_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacccccccc)
  ) CLBLM_R_X27Y14_SLICE_X43Y14_CLUT (
.I0(CLBLM_R_X27Y14_SLICE_X43Y14_AQ),
.I1(CLBLM_R_X27Y14_SLICE_X43Y14_B_XOR),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y14_SLICE_X43Y14_CO5),
.O6(CLBLM_R_X27Y14_SLICE_X43Y14_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X27Y14_SLICE_X43Y14_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y14_SLICE_X43Y14_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y14_SLICE_X43Y14_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X27Y14_SLICE_X43Y14_BO5),
.O6(CLBLM_R_X27Y14_SLICE_X43Y14_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0fffff0000)
  ) CLBLM_R_X27Y14_SLICE_X43Y14_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X27Y14_SLICE_X43Y14_DQ),
.I3(1'b1),
.I4(CLBLM_R_X27Y14_SLICE_X43Y14_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X27Y14_SLICE_X43Y14_AO5),
.O6(CLBLM_R_X27Y14_SLICE_X43Y14_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y15_SLICE_X42Y15_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y15_SLICE_X42Y15_DO5),
.O6(CLBLM_R_X27Y15_SLICE_X42Y15_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y15_SLICE_X42Y15_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y15_SLICE_X42Y15_CO5),
.O6(CLBLM_R_X27Y15_SLICE_X42Y15_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y15_SLICE_X42Y15_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y15_SLICE_X42Y15_BO5),
.O6(CLBLM_R_X27Y15_SLICE_X42Y15_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y15_SLICE_X42Y15_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y15_SLICE_X42Y15_AO5),
.O6(CLBLM_R_X27Y15_SLICE_X42Y15_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y15_SLICE_X43Y15_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y15_SLICE_X43Y15_AO5),
.Q(CLBLM_R_X27Y15_SLICE_X43Y15_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y15_SLICE_X43Y15_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y15_SLICE_X43Y15_BO5),
.Q(CLBLM_R_X27Y15_SLICE_X43Y15_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y15_SLICE_X43Y15_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y15_SLICE_X43Y15_CO5),
.Q(CLBLM_R_X27Y15_SLICE_X43Y15_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y15_SLICE_X43Y15_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y15_SLICE_X43Y15_DO5),
.Q(CLBLM_R_X27Y15_SLICE_X43Y15_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X27Y15_SLICE_X43Y15_CARRY4 (
.CI(CLBLM_R_X27Y14_SLICE_X43Y14_COUT),
.CO({CLBLM_R_X27Y15_SLICE_X43Y15_D_CY, CLBLM_R_X27Y15_SLICE_X43Y15_C_CY, CLBLM_R_X27Y15_SLICE_X43Y15_B_CY, CLBLM_R_X27Y15_SLICE_X43Y15_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X27Y15_SLICE_X43Y15_D_XOR, CLBLM_R_X27Y15_SLICE_X43Y15_C_XOR, CLBLM_R_X27Y15_SLICE_X43Y15_B_XOR, CLBLM_R_X27Y15_SLICE_X43Y15_A_XOR}),
.S({CLBLM_R_X27Y15_SLICE_X43Y15_DO6, CLBLM_R_X27Y15_SLICE_X43Y15_CO6, CLBLM_R_X27Y15_SLICE_X43Y15_BO6, CLBLM_R_X27Y15_SLICE_X43Y15_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLM_R_X27Y15_SLICE_X43Y15_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X27Y15_SLICE_X43Y15_B_XOR),
.I4(CLBLM_R_X27Y15_SLICE_X43Y15_BQ),
.I5(1'b1),
.O5(CLBLM_R_X27Y15_SLICE_X43Y15_DO5),
.O6(CLBLM_R_X27Y15_SLICE_X43Y15_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X27Y15_SLICE_X43Y15_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y15_SLICE_X43Y15_A_XOR),
.I2(CLBLM_R_X27Y15_SLICE_X43Y15_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y15_SLICE_X43Y15_CO5),
.O6(CLBLM_R_X27Y15_SLICE_X43Y15_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X27Y15_SLICE_X43Y15_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y15_SLICE_X43Y15_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y15_SLICE_X43Y15_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X27Y15_SLICE_X43Y15_BO5),
.O6(CLBLM_R_X27Y15_SLICE_X43Y15_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X27Y15_SLICE_X43Y15_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y15_SLICE_X43Y15_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y15_SLICE_X43Y15_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X27Y15_SLICE_X43Y15_AO5),
.O6(CLBLM_R_X27Y15_SLICE_X43Y15_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y16_SLICE_X42Y16_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y16_SLICE_X42Y16_DO5),
.O6(CLBLM_R_X27Y16_SLICE_X42Y16_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y16_SLICE_X42Y16_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y16_SLICE_X42Y16_CO5),
.O6(CLBLM_R_X27Y16_SLICE_X42Y16_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y16_SLICE_X42Y16_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y16_SLICE_X42Y16_BO5),
.O6(CLBLM_R_X27Y16_SLICE_X42Y16_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y16_SLICE_X42Y16_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y16_SLICE_X42Y16_AO5),
.O6(CLBLM_R_X27Y16_SLICE_X42Y16_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y16_SLICE_X43Y16_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y16_SLICE_X43Y16_AO5),
.Q(CLBLM_R_X27Y16_SLICE_X43Y16_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y16_SLICE_X43Y16_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y16_SLICE_X43Y16_BO5),
.Q(CLBLM_R_X27Y16_SLICE_X43Y16_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y16_SLICE_X43Y16_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y16_SLICE_X43Y16_CO5),
.Q(CLBLM_R_X27Y16_SLICE_X43Y16_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y16_SLICE_X43Y16_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y16_SLICE_X43Y16_DO5),
.Q(CLBLM_R_X27Y16_SLICE_X43Y16_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X27Y16_SLICE_X43Y16_CARRY4 (
.CI(CLBLM_R_X27Y15_SLICE_X43Y15_COUT),
.CO({CLBLM_R_X27Y16_SLICE_X43Y16_D_CY, CLBLM_R_X27Y16_SLICE_X43Y16_C_CY, CLBLM_R_X27Y16_SLICE_X43Y16_B_CY, CLBLM_R_X27Y16_SLICE_X43Y16_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X27Y16_SLICE_X43Y16_D_XOR, CLBLM_R_X27Y16_SLICE_X43Y16_C_XOR, CLBLM_R_X27Y16_SLICE_X43Y16_B_XOR, CLBLM_R_X27Y16_SLICE_X43Y16_A_XOR}),
.S({CLBLM_R_X27Y16_SLICE_X43Y16_DO6, CLBLM_R_X27Y16_SLICE_X43Y16_CO6, CLBLM_R_X27Y16_SLICE_X43Y16_BO6, CLBLM_R_X27Y16_SLICE_X43Y16_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLM_R_X27Y16_SLICE_X43Y16_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X27Y16_SLICE_X43Y16_B_XOR),
.I4(CLBLM_R_X27Y16_SLICE_X43Y16_BQ),
.I5(1'b1),
.O5(CLBLM_R_X27Y16_SLICE_X43Y16_DO5),
.O6(CLBLM_R_X27Y16_SLICE_X43Y16_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X27Y16_SLICE_X43Y16_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y16_SLICE_X43Y16_A_XOR),
.I2(CLBLM_R_X27Y16_SLICE_X43Y16_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y16_SLICE_X43Y16_CO5),
.O6(CLBLM_R_X27Y16_SLICE_X43Y16_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X27Y16_SLICE_X43Y16_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y16_SLICE_X43Y16_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y16_SLICE_X43Y16_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X27Y16_SLICE_X43Y16_BO5),
.O6(CLBLM_R_X27Y16_SLICE_X43Y16_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X27Y16_SLICE_X43Y16_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y16_SLICE_X43Y16_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y16_SLICE_X43Y16_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X27Y16_SLICE_X43Y16_AO5),
.O6(CLBLM_R_X27Y16_SLICE_X43Y16_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y17_SLICE_X42Y17_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y17_SLICE_X42Y17_DO5),
.O6(CLBLM_R_X27Y17_SLICE_X42Y17_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y17_SLICE_X42Y17_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y17_SLICE_X42Y17_CO5),
.O6(CLBLM_R_X27Y17_SLICE_X42Y17_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y17_SLICE_X42Y17_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y17_SLICE_X42Y17_BO5),
.O6(CLBLM_R_X27Y17_SLICE_X42Y17_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y17_SLICE_X42Y17_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y17_SLICE_X42Y17_AO5),
.O6(CLBLM_R_X27Y17_SLICE_X42Y17_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y17_SLICE_X43Y17_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y17_SLICE_X43Y17_A_XOR),
.Q(CLBLM_R_X27Y17_SLICE_X43Y17_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y17_SLICE_X43Y17_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y17_SLICE_X43Y17_BO5),
.Q(CLBLM_R_X27Y17_SLICE_X43Y17_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y17_SLICE_X43Y17_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y17_SLICE_X43Y17_CO5),
.Q(CLBLM_R_X27Y17_SLICE_X43Y17_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y17_SLICE_X43Y17_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y17_SLICE_X43Y17_DO5),
.Q(CLBLM_R_X27Y17_SLICE_X43Y17_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X27Y17_SLICE_X43Y17_CARRY4 (
.CI(CLBLM_R_X27Y16_SLICE_X43Y16_COUT),
.CO({CLBLM_R_X27Y17_SLICE_X43Y17_D_CY, CLBLM_R_X27Y17_SLICE_X43Y17_C_CY, CLBLM_R_X27Y17_SLICE_X43Y17_B_CY, CLBLM_R_X27Y17_SLICE_X43Y17_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X27Y17_SLICE_X43Y17_D_XOR, CLBLM_R_X27Y17_SLICE_X43Y17_C_XOR, CLBLM_R_X27Y17_SLICE_X43Y17_B_XOR, CLBLM_R_X27Y17_SLICE_X43Y17_A_XOR}),
.S({CLBLM_R_X27Y17_SLICE_X43Y17_DO6, CLBLM_R_X27Y17_SLICE_X43Y17_CO6, CLBLM_R_X27Y17_SLICE_X43Y17_BO6, CLBLM_R_X27Y17_SLICE_X43Y17_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X27Y17_SLICE_X43Y17_DLUT (
.I0(CLBLM_R_X27Y17_SLICE_X43Y17_B_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y17_SLICE_X43Y17_CQ),
.I5(1'b1),
.O5(CLBLM_R_X27Y17_SLICE_X43Y17_DO5),
.O6(CLBLM_R_X27Y17_SLICE_X43Y17_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X27Y17_SLICE_X43Y17_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y17_SLICE_X43Y17_D_XOR),
.I2(CLBLM_R_X27Y17_SLICE_X43Y17_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y17_SLICE_X43Y17_CO5),
.O6(CLBLM_R_X27Y17_SLICE_X43Y17_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLM_R_X27Y17_SLICE_X43Y17_BLUT (
.I0(CLBLM_R_X27Y17_SLICE_X43Y17_C_XOR),
.I1(CLBLM_R_X27Y17_SLICE_X43Y17_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y17_SLICE_X43Y17_BO5),
.O6(CLBLM_R_X27Y17_SLICE_X43Y17_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X27Y17_SLICE_X43Y17_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y17_SLICE_X43Y17_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y17_SLICE_X43Y17_AO5),
.O6(CLBLM_R_X27Y17_SLICE_X43Y17_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y18_SLICE_X42Y18_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y18_SLICE_X42Y18_DO5),
.O6(CLBLM_R_X27Y18_SLICE_X42Y18_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y18_SLICE_X42Y18_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y18_SLICE_X42Y18_CO5),
.O6(CLBLM_R_X27Y18_SLICE_X42Y18_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y18_SLICE_X42Y18_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y18_SLICE_X42Y18_BO5),
.O6(CLBLM_R_X27Y18_SLICE_X42Y18_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y18_SLICE_X42Y18_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y18_SLICE_X42Y18_AO5),
.O6(CLBLM_R_X27Y18_SLICE_X42Y18_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y18_SLICE_X43Y18_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y18_SLICE_X43Y18_A_XOR),
.Q(CLBLM_R_X27Y18_SLICE_X43Y18_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y18_SLICE_X43Y18_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y18_SLICE_X43Y18_BO5),
.Q(CLBLM_R_X27Y18_SLICE_X43Y18_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y18_SLICE_X43Y18_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y18_SLICE_X43Y18_CO5),
.Q(CLBLM_R_X27Y18_SLICE_X43Y18_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y18_SLICE_X43Y18_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y18_SLICE_X43Y18_DO5),
.Q(CLBLM_R_X27Y18_SLICE_X43Y18_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X27Y18_SLICE_X43Y18_CARRY4 (
.CI(CLBLM_R_X27Y17_SLICE_X43Y17_COUT),
.CO({CLBLM_R_X27Y18_SLICE_X43Y18_D_CY, CLBLM_R_X27Y18_SLICE_X43Y18_C_CY, CLBLM_R_X27Y18_SLICE_X43Y18_B_CY, CLBLM_R_X27Y18_SLICE_X43Y18_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X27Y18_SLICE_X43Y18_D_XOR, CLBLM_R_X27Y18_SLICE_X43Y18_C_XOR, CLBLM_R_X27Y18_SLICE_X43Y18_B_XOR, CLBLM_R_X27Y18_SLICE_X43Y18_A_XOR}),
.S({CLBLM_R_X27Y18_SLICE_X43Y18_DO6, CLBLM_R_X27Y18_SLICE_X43Y18_CO6, CLBLM_R_X27Y18_SLICE_X43Y18_BO6, CLBLM_R_X27Y18_SLICE_X43Y18_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X27Y18_SLICE_X43Y18_DLUT (
.I0(CLBLM_R_X27Y18_SLICE_X43Y18_B_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y18_SLICE_X43Y18_CQ),
.I5(1'b1),
.O5(CLBLM_R_X27Y18_SLICE_X43Y18_DO5),
.O6(CLBLM_R_X27Y18_SLICE_X43Y18_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X27Y18_SLICE_X43Y18_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y18_SLICE_X43Y18_D_XOR),
.I2(CLBLM_R_X27Y18_SLICE_X43Y18_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y18_SLICE_X43Y18_CO5),
.O6(CLBLM_R_X27Y18_SLICE_X43Y18_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLM_R_X27Y18_SLICE_X43Y18_BLUT (
.I0(CLBLM_R_X27Y18_SLICE_X43Y18_C_XOR),
.I1(CLBLM_R_X27Y18_SLICE_X43Y18_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y18_SLICE_X43Y18_BO5),
.O6(CLBLM_R_X27Y18_SLICE_X43Y18_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X27Y18_SLICE_X43Y18_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y18_SLICE_X43Y18_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y18_SLICE_X43Y18_AO5),
.O6(CLBLM_R_X27Y18_SLICE_X43Y18_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y19_SLICE_X42Y19_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y19_SLICE_X42Y19_DO5),
.O6(CLBLM_R_X27Y19_SLICE_X42Y19_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y19_SLICE_X42Y19_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y19_SLICE_X42Y19_CO5),
.O6(CLBLM_R_X27Y19_SLICE_X42Y19_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y19_SLICE_X42Y19_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y19_SLICE_X42Y19_BO5),
.O6(CLBLM_R_X27Y19_SLICE_X42Y19_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y19_SLICE_X42Y19_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y19_SLICE_X42Y19_AO5),
.O6(CLBLM_R_X27Y19_SLICE_X42Y19_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y19_SLICE_X43Y19_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y19_SLICE_X43Y19_AO5),
.Q(CLBLM_R_X27Y19_SLICE_X43Y19_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y19_SLICE_X43Y19_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y19_SLICE_X43Y19_BO5),
.Q(CLBLM_R_X27Y19_SLICE_X43Y19_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y19_SLICE_X43Y19_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y19_SLICE_X43Y19_C_XOR),
.Q(CLBLM_R_X27Y19_SLICE_X43Y19_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y19_SLICE_X43Y19_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y19_SLICE_X43Y19_D_XOR),
.Q(CLBLM_R_X27Y19_SLICE_X43Y19_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X27Y19_SLICE_X43Y19_CARRY4 (
.CI(CLBLM_R_X27Y18_SLICE_X43Y18_COUT),
.CO({CLBLM_R_X27Y19_SLICE_X43Y19_D_CY, CLBLM_R_X27Y19_SLICE_X43Y19_C_CY, CLBLM_R_X27Y19_SLICE_X43Y19_B_CY, CLBLM_R_X27Y19_SLICE_X43Y19_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X27Y19_SLICE_X43Y19_D_XOR, CLBLM_R_X27Y19_SLICE_X43Y19_C_XOR, CLBLM_R_X27Y19_SLICE_X43Y19_B_XOR, CLBLM_R_X27Y19_SLICE_X43Y19_A_XOR}),
.S({CLBLM_R_X27Y19_SLICE_X43Y19_DO6, CLBLM_R_X27Y19_SLICE_X43Y19_CO6, CLBLM_R_X27Y19_SLICE_X43Y19_BO6, CLBLM_R_X27Y19_SLICE_X43Y19_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff000000000000)
  ) CLBLM_R_X27Y19_SLICE_X43Y19_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y19_SLICE_X43Y19_DQ),
.I5(1'b1),
.O5(CLBLM_R_X27Y19_SLICE_X43Y19_DO5),
.O6(CLBLM_R_X27Y19_SLICE_X43Y19_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ccccffff)
  ) CLBLM_R_X27Y19_SLICE_X43Y19_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y8_SLICE_X42Y8_DQ),
.I2(CLBLM_R_X27Y19_SLICE_X43Y19_CQ),
.I3(1'b1),
.I4(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_LOCKED),
.I5(1'b1),
.O5(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.O6(CLBLM_R_X27Y19_SLICE_X43Y19_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X27Y19_SLICE_X43Y19_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y19_SLICE_X43Y19_AQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y19_SLICE_X43Y19_A_XOR),
.I5(1'b1),
.O5(CLBLM_R_X27Y19_SLICE_X43Y19_BO5),
.O6(CLBLM_R_X27Y19_SLICE_X43Y19_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X27Y19_SLICE_X43Y19_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y19_SLICE_X43Y19_BQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y19_SLICE_X43Y19_B_XOR),
.I5(1'b1),
.O5(CLBLM_R_X27Y19_SLICE_X43Y19_AO5),
.O6(CLBLM_R_X27Y19_SLICE_X43Y19_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y38_SLICE_X42Y38_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y38_SLICE_X42Y38_DO5),
.O6(CLBLM_R_X27Y38_SLICE_X42Y38_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y38_SLICE_X42Y38_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y38_SLICE_X42Y38_CO5),
.O6(CLBLM_R_X27Y38_SLICE_X42Y38_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y38_SLICE_X42Y38_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y38_SLICE_X42Y38_BO5),
.O6(CLBLM_R_X27Y38_SLICE_X42Y38_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y38_SLICE_X42Y38_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y38_SLICE_X42Y38_AO5),
.O6(CLBLM_R_X27Y38_SLICE_X42Y38_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y38_SLICE_X43Y38_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y38_SLICE_X43Y38_AO5),
.Q(CLBLM_R_X27Y38_SLICE_X43Y38_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y38_SLICE_X43Y38_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y38_SLICE_X43Y38_BO5),
.Q(CLBLM_R_X27Y38_SLICE_X43Y38_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y38_SLICE_X43Y38_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y38_SLICE_X43Y38_CO5),
.Q(CLBLM_R_X27Y38_SLICE_X43Y38_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y38_SLICE_X43Y38_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y38_SLICE_X43Y38_DO5),
.Q(CLBLM_R_X27Y38_SLICE_X43Y38_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X27Y38_SLICE_X43Y38_CARRY4 (
.CI(1'b0),
.CO({CLBLM_R_X27Y38_SLICE_X43Y38_D_CY, CLBLM_R_X27Y38_SLICE_X43Y38_C_CY, CLBLM_R_X27Y38_SLICE_X43Y38_B_CY, CLBLM_R_X27Y38_SLICE_X43Y38_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b1}),
.O({CLBLM_R_X27Y38_SLICE_X43Y38_D_XOR, CLBLM_R_X27Y38_SLICE_X43Y38_C_XOR, CLBLM_R_X27Y38_SLICE_X43Y38_B_XOR, CLBLM_R_X27Y38_SLICE_X43Y38_A_XOR}),
.S({CLBLM_R_X27Y38_SLICE_X43Y38_DO6, CLBLM_R_X27Y38_SLICE_X43Y38_CO6, CLBLM_R_X27Y38_SLICE_X43Y38_BO6, CLBLM_R_X27Y38_SLICE_X43Y38_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X27Y38_SLICE_X43Y38_DLUT (
.I0(CLBLM_R_X27Y38_SLICE_X43Y38_AO6),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y38_SLICE_X43Y38_CQ),
.I5(1'b1),
.O5(CLBLM_R_X27Y38_SLICE_X43Y38_DO5),
.O6(CLBLM_R_X27Y38_SLICE_X43Y38_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'haaaaaaaacccccccc)
  ) CLBLM_R_X27Y38_SLICE_X43Y38_CLUT (
.I0(CLBLM_R_X27Y42_SLICE_X43Y42_A5Q),
.I1(CLBLM_R_X27Y38_SLICE_X43Y38_D_XOR),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y38_SLICE_X43Y38_CO5),
.O6(CLBLM_R_X27Y38_SLICE_X43Y38_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0ff00ff00)
  ) CLBLM_R_X27Y38_SLICE_X43Y38_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLM_R_X27Y41_SLICE_X43Y41_A5Q),
.I3(CLBLM_R_X27Y43_SLICE_X43Y43_D_XOR),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y38_SLICE_X43Y38_BO5),
.O6(CLBLM_R_X27Y38_SLICE_X43Y38_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0f0f0faaaaaaaa)
  ) CLBLM_R_X27Y38_SLICE_X43Y38_ALUT (
.I0(CLBLM_R_X27Y43_SLICE_X43Y43_C_XOR),
.I1(1'b1),
.I2(CLBLM_R_X27Y38_SLICE_X43Y38_DQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y38_SLICE_X43Y38_AO5),
.O6(CLBLM_R_X27Y38_SLICE_X43Y38_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y39_SLICE_X42Y39_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y39_SLICE_X42Y39_DO5),
.O6(CLBLM_R_X27Y39_SLICE_X42Y39_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y39_SLICE_X42Y39_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y39_SLICE_X42Y39_CO5),
.O6(CLBLM_R_X27Y39_SLICE_X42Y39_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y39_SLICE_X42Y39_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y39_SLICE_X42Y39_BO5),
.O6(CLBLM_R_X27Y39_SLICE_X42Y39_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y39_SLICE_X42Y39_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y39_SLICE_X42Y39_AO5),
.O6(CLBLM_R_X27Y39_SLICE_X42Y39_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y39_SLICE_X43Y39_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y39_SLICE_X43Y39_AO5),
.Q(CLBLM_R_X27Y39_SLICE_X43Y39_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y39_SLICE_X43Y39_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y39_SLICE_X43Y39_BO5),
.Q(CLBLM_R_X27Y39_SLICE_X43Y39_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y39_SLICE_X43Y39_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y39_SLICE_X43Y39_CO5),
.Q(CLBLM_R_X27Y39_SLICE_X43Y39_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y39_SLICE_X43Y39_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y39_SLICE_X43Y39_DO5),
.Q(CLBLM_R_X27Y39_SLICE_X43Y39_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X27Y39_SLICE_X43Y39_CARRY4 (
.CI(CLBLM_R_X27Y38_SLICE_X43Y38_COUT),
.CO({CLBLM_R_X27Y39_SLICE_X43Y39_D_CY, CLBLM_R_X27Y39_SLICE_X43Y39_C_CY, CLBLM_R_X27Y39_SLICE_X43Y39_B_CY, CLBLM_R_X27Y39_SLICE_X43Y39_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X27Y39_SLICE_X43Y39_D_XOR, CLBLM_R_X27Y39_SLICE_X43Y39_C_XOR, CLBLM_R_X27Y39_SLICE_X43Y39_B_XOR, CLBLM_R_X27Y39_SLICE_X43Y39_A_XOR}),
.S({CLBLM_R_X27Y39_SLICE_X43Y39_DO6, CLBLM_R_X27Y39_SLICE_X43Y39_CO6, CLBLM_R_X27Y39_SLICE_X43Y39_BO6, CLBLM_R_X27Y39_SLICE_X43Y39_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLM_R_X27Y39_SLICE_X43Y39_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X27Y39_SLICE_X43Y39_B_XOR),
.I4(CLBLM_R_X27Y39_SLICE_X43Y39_BQ),
.I5(1'b1),
.O5(CLBLM_R_X27Y39_SLICE_X43Y39_DO5),
.O6(CLBLM_R_X27Y39_SLICE_X43Y39_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X27Y39_SLICE_X43Y39_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y39_SLICE_X43Y39_A_XOR),
.I2(CLBLM_R_X27Y39_SLICE_X43Y39_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y39_SLICE_X43Y39_CO5),
.O6(CLBLM_R_X27Y39_SLICE_X43Y39_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X27Y39_SLICE_X43Y39_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y39_SLICE_X43Y39_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y39_SLICE_X43Y39_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X27Y39_SLICE_X43Y39_BO5),
.O6(CLBLM_R_X27Y39_SLICE_X43Y39_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X27Y39_SLICE_X43Y39_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y39_SLICE_X43Y39_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y39_SLICE_X43Y39_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X27Y39_SLICE_X43Y39_AO5),
.O6(CLBLM_R_X27Y39_SLICE_X43Y39_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y40_SLICE_X42Y40_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y40_SLICE_X42Y40_DO5),
.O6(CLBLM_R_X27Y40_SLICE_X42Y40_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y40_SLICE_X42Y40_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y40_SLICE_X42Y40_CO5),
.O6(CLBLM_R_X27Y40_SLICE_X42Y40_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y40_SLICE_X42Y40_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y40_SLICE_X42Y40_BO5),
.O6(CLBLM_R_X27Y40_SLICE_X42Y40_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y40_SLICE_X42Y40_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y40_SLICE_X42Y40_AO5),
.O6(CLBLM_R_X27Y40_SLICE_X42Y40_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y40_SLICE_X43Y40_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y40_SLICE_X43Y40_AO5),
.Q(CLBLM_R_X27Y40_SLICE_X43Y40_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y40_SLICE_X43Y40_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y40_SLICE_X43Y40_BO5),
.Q(CLBLM_R_X27Y40_SLICE_X43Y40_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y40_SLICE_X43Y40_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y40_SLICE_X43Y40_CO5),
.Q(CLBLM_R_X27Y40_SLICE_X43Y40_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y40_SLICE_X43Y40_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y40_SLICE_X43Y40_DO5),
.Q(CLBLM_R_X27Y40_SLICE_X43Y40_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X27Y40_SLICE_X43Y40_CARRY4 (
.CI(CLBLM_R_X27Y39_SLICE_X43Y39_COUT),
.CO({CLBLM_R_X27Y40_SLICE_X43Y40_D_CY, CLBLM_R_X27Y40_SLICE_X43Y40_C_CY, CLBLM_R_X27Y40_SLICE_X43Y40_B_CY, CLBLM_R_X27Y40_SLICE_X43Y40_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X27Y40_SLICE_X43Y40_D_XOR, CLBLM_R_X27Y40_SLICE_X43Y40_C_XOR, CLBLM_R_X27Y40_SLICE_X43Y40_B_XOR, CLBLM_R_X27Y40_SLICE_X43Y40_A_XOR}),
.S({CLBLM_R_X27Y40_SLICE_X43Y40_DO6, CLBLM_R_X27Y40_SLICE_X43Y40_CO6, CLBLM_R_X27Y40_SLICE_X43Y40_BO6, CLBLM_R_X27Y40_SLICE_X43Y40_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLM_R_X27Y40_SLICE_X43Y40_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X27Y40_SLICE_X43Y40_B_XOR),
.I4(CLBLM_R_X27Y40_SLICE_X43Y40_BQ),
.I5(1'b1),
.O5(CLBLM_R_X27Y40_SLICE_X43Y40_DO5),
.O6(CLBLM_R_X27Y40_SLICE_X43Y40_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X27Y40_SLICE_X43Y40_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y40_SLICE_X43Y40_A_XOR),
.I2(CLBLM_R_X27Y40_SLICE_X43Y40_AQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y40_SLICE_X43Y40_CO5),
.O6(CLBLM_R_X27Y40_SLICE_X43Y40_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X27Y40_SLICE_X43Y40_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y40_SLICE_X43Y40_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y40_SLICE_X43Y40_D_XOR),
.I5(1'b1),
.O5(CLBLM_R_X27Y40_SLICE_X43Y40_BO5),
.O6(CLBLM_R_X27Y40_SLICE_X43Y40_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccffff0000)
  ) CLBLM_R_X27Y40_SLICE_X43Y40_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y40_SLICE_X43Y40_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y40_SLICE_X43Y40_C_XOR),
.I5(1'b1),
.O5(CLBLM_R_X27Y40_SLICE_X43Y40_AO5),
.O6(CLBLM_R_X27Y40_SLICE_X43Y40_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y41_SLICE_X42Y41_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y41_SLICE_X42Y41_DO5),
.O6(CLBLM_R_X27Y41_SLICE_X42Y41_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y41_SLICE_X42Y41_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y41_SLICE_X42Y41_CO5),
.O6(CLBLM_R_X27Y41_SLICE_X42Y41_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y41_SLICE_X42Y41_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y41_SLICE_X42Y41_BO5),
.O6(CLBLM_R_X27Y41_SLICE_X42Y41_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y41_SLICE_X42Y41_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y41_SLICE_X42Y41_AO5),
.O6(CLBLM_R_X27Y41_SLICE_X42Y41_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y41_SLICE_X43Y41_A5_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y41_SLICE_X43Y41_AO5),
.Q(CLBLM_R_X27Y41_SLICE_X43Y41_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y41_SLICE_X43Y41_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y41_SLICE_X43Y41_A_XOR),
.Q(CLBLM_R_X27Y41_SLICE_X43Y41_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y41_SLICE_X43Y41_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y41_SLICE_X43Y41_BO5),
.Q(CLBLM_R_X27Y41_SLICE_X43Y41_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y41_SLICE_X43Y41_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y41_SLICE_X43Y41_CO5),
.Q(CLBLM_R_X27Y41_SLICE_X43Y41_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y41_SLICE_X43Y41_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y41_SLICE_X43Y41_DO5),
.Q(CLBLM_R_X27Y41_SLICE_X43Y41_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X27Y41_SLICE_X43Y41_CARRY4 (
.CI(CLBLM_R_X27Y40_SLICE_X43Y40_COUT),
.CO({CLBLM_R_X27Y41_SLICE_X43Y41_D_CY, CLBLM_R_X27Y41_SLICE_X43Y41_C_CY, CLBLM_R_X27Y41_SLICE_X43Y41_B_CY, CLBLM_R_X27Y41_SLICE_X43Y41_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X27Y41_SLICE_X43Y41_D_XOR, CLBLM_R_X27Y41_SLICE_X43Y41_C_XOR, CLBLM_R_X27Y41_SLICE_X43Y41_B_XOR, CLBLM_R_X27Y41_SLICE_X43Y41_A_XOR}),
.S({CLBLM_R_X27Y41_SLICE_X43Y41_DO6, CLBLM_R_X27Y41_SLICE_X43Y41_CO6, CLBLM_R_X27Y41_SLICE_X43Y41_BO6, CLBLM_R_X27Y41_SLICE_X43Y41_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X27Y41_SLICE_X43Y41_DLUT (
.I0(CLBLM_R_X27Y41_SLICE_X43Y41_B_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y41_SLICE_X43Y41_CQ),
.I5(1'b1),
.O5(CLBLM_R_X27Y41_SLICE_X43Y41_DO5),
.O6(CLBLM_R_X27Y41_SLICE_X43Y41_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X27Y41_SLICE_X43Y41_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y41_SLICE_X43Y41_D_XOR),
.I2(CLBLM_R_X27Y41_SLICE_X43Y41_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y41_SLICE_X43Y41_CO5),
.O6(CLBLM_R_X27Y41_SLICE_X43Y41_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLM_R_X27Y41_SLICE_X43Y41_BLUT (
.I0(CLBLM_R_X27Y41_SLICE_X43Y41_C_XOR),
.I1(CLBLM_R_X27Y41_SLICE_X43Y41_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y41_SLICE_X43Y41_BO5),
.O6(CLBLM_R_X27Y41_SLICE_X43Y41_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0f0f0f0)
  ) CLBLM_R_X27Y41_SLICE_X43Y41_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y41_SLICE_X43Y41_AQ),
.I2(CLBLM_R_X27Y38_SLICE_X43Y38_B_XOR),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y41_SLICE_X43Y41_AO5),
.O6(CLBLM_R_X27Y41_SLICE_X43Y41_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y42_SLICE_X42Y42_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y42_SLICE_X42Y42_DO5),
.O6(CLBLM_R_X27Y42_SLICE_X42Y42_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y42_SLICE_X42Y42_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y42_SLICE_X42Y42_CO5),
.O6(CLBLM_R_X27Y42_SLICE_X42Y42_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y42_SLICE_X42Y42_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y42_SLICE_X42Y42_BO5),
.O6(CLBLM_R_X27Y42_SLICE_X42Y42_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y42_SLICE_X42Y42_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y42_SLICE_X42Y42_AO5),
.O6(CLBLM_R_X27Y42_SLICE_X42Y42_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A5FF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y42_SLICE_X43Y42_A5_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y42_SLICE_X43Y42_AO5),
.Q(CLBLM_R_X27Y42_SLICE_X43Y42_A5Q)
  );


  (* KEEP, DONT_TOUCH, BEL = "AFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y42_SLICE_X43Y42_A_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y42_SLICE_X43Y42_A_XOR),
.Q(CLBLM_R_X27Y42_SLICE_X43Y42_AQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "BFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y42_SLICE_X43Y42_B_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y42_SLICE_X43Y42_BO5),
.Q(CLBLM_R_X27Y42_SLICE_X43Y42_BQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y42_SLICE_X43Y42_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y42_SLICE_X43Y42_CO5),
.Q(CLBLM_R_X27Y42_SLICE_X43Y42_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y42_SLICE_X43Y42_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y42_SLICE_X43Y42_DO5),
.Q(CLBLM_R_X27Y42_SLICE_X43Y42_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X27Y42_SLICE_X43Y42_CARRY4 (
.CI(CLBLM_R_X27Y41_SLICE_X43Y41_COUT),
.CO({CLBLM_R_X27Y42_SLICE_X43Y42_D_CY, CLBLM_R_X27Y42_SLICE_X43Y42_C_CY, CLBLM_R_X27Y42_SLICE_X43Y42_B_CY, CLBLM_R_X27Y42_SLICE_X43Y42_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X27Y42_SLICE_X43Y42_D_XOR, CLBLM_R_X27Y42_SLICE_X43Y42_C_XOR, CLBLM_R_X27Y42_SLICE_X43Y42_B_XOR, CLBLM_R_X27Y42_SLICE_X43Y42_A_XOR}),
.S({CLBLM_R_X27Y42_SLICE_X43Y42_DO6, CLBLM_R_X27Y42_SLICE_X43Y42_CO6, CLBLM_R_X27Y42_SLICE_X43Y42_BO6, CLBLM_R_X27Y42_SLICE_X43Y42_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000aaaaaaaa)
  ) CLBLM_R_X27Y42_SLICE_X43Y42_DLUT (
.I0(CLBLM_R_X27Y42_SLICE_X43Y42_B_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(CLBLM_R_X27Y42_SLICE_X43Y42_CQ),
.I5(1'b1),
.O5(CLBLM_R_X27Y42_SLICE_X43Y42_DO5),
.O6(CLBLM_R_X27Y42_SLICE_X43Y42_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f0f0f0cccccccc)
  ) CLBLM_R_X27Y42_SLICE_X43Y42_CLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y42_SLICE_X43Y42_D_XOR),
.I2(CLBLM_R_X27Y42_SLICE_X43Y42_BQ),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y42_SLICE_X43Y42_CO5),
.O6(CLBLM_R_X27Y42_SLICE_X43Y42_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccaaaaaaaa)
  ) CLBLM_R_X27Y42_SLICE_X43Y42_BLUT (
.I0(CLBLM_R_X27Y42_SLICE_X43Y42_C_XOR),
.I1(CLBLM_R_X27Y42_SLICE_X43Y42_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y42_SLICE_X43Y42_BO5),
.O6(CLBLM_R_X27Y42_SLICE_X43Y42_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hccccccccf0f0f0f0)
  ) CLBLM_R_X27Y42_SLICE_X43Y42_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y42_SLICE_X43Y42_AQ),
.I2(CLBLM_R_X27Y38_SLICE_X43Y38_C_XOR),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y42_SLICE_X43Y42_AO5),
.O6(CLBLM_R_X27Y42_SLICE_X43Y42_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y43_SLICE_X42Y43_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y43_SLICE_X42Y43_DO5),
.O6(CLBLM_R_X27Y43_SLICE_X42Y43_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y43_SLICE_X42Y43_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y43_SLICE_X42Y43_CO5),
.O6(CLBLM_R_X27Y43_SLICE_X42Y43_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y43_SLICE_X42Y43_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y43_SLICE_X42Y43_BO5),
.O6(CLBLM_R_X27Y43_SLICE_X42Y43_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLM_R_X27Y43_SLICE_X42Y43_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y43_SLICE_X42Y43_AO5),
.O6(CLBLM_R_X27Y43_SLICE_X42Y43_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "CFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y43_SLICE_X43Y43_C_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y43_SLICE_X43Y43_CO5),
.Q(CLBLM_R_X27Y43_SLICE_X43Y43_CQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "DFF" *)
  FDCE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLM_R_X27Y43_SLICE_X43Y43_D_FDCE (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O),
.CE(1'b1),
.CLR(CLBLM_R_X27Y19_SLICE_X43Y19_CO5),
.D(CLBLM_R_X27Y43_SLICE_X43Y43_DO5),
.Q(CLBLM_R_X27Y43_SLICE_X43Y43_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLM_R_X27Y43_SLICE_X43Y43_CARRY4 (
.CI(CLBLM_R_X27Y42_SLICE_X43Y42_COUT),
.CO({CLBLM_R_X27Y43_SLICE_X43Y43_D_CY, CLBLM_R_X27Y43_SLICE_X43Y43_C_CY, CLBLM_R_X27Y43_SLICE_X43Y43_B_CY, CLBLM_R_X27Y43_SLICE_X43Y43_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0}),
.O({CLBLM_R_X27Y43_SLICE_X43Y43_D_XOR, CLBLM_R_X27Y43_SLICE_X43Y43_C_XOR, CLBLM_R_X27Y43_SLICE_X43Y43_B_XOR, CLBLM_R_X27Y43_SLICE_X43Y43_A_XOR}),
.S({CLBLM_R_X27Y43_SLICE_X43Y43_DO6, CLBLM_R_X27Y43_SLICE_X43Y43_CO6, CLBLM_R_X27Y43_SLICE_X43Y43_BO6, CLBLM_R_X27Y43_SLICE_X43Y43_AO6})
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'hffff0000ff00ff00)
  ) CLBLM_R_X27Y43_SLICE_X43Y43_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X27Y43_SLICE_X43Y43_A_XOR),
.I4(CLBLM_R_X27Y38_SLICE_X43Y38_BQ),
.I5(1'b1),
.O5(CLBLM_R_X27Y43_SLICE_X43Y43_DO5),
.O6(CLBLM_R_X27Y43_SLICE_X43Y43_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'hff00ff00aaaaaaaa)
  ) CLBLM_R_X27Y43_SLICE_X43Y43_CLUT (
.I0(CLBLM_R_X27Y43_SLICE_X43Y43_B_XOR),
.I1(1'b1),
.I2(1'b1),
.I3(CLBLM_R_X27Y38_SLICE_X43Y38_AQ),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y43_SLICE_X43Y43_CO5),
.O6(CLBLM_R_X27Y43_SLICE_X43Y43_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X27Y43_SLICE_X43Y43_BLUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y43_SLICE_X43Y43_CQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y43_SLICE_X43Y43_BO5),
.O6(CLBLM_R_X27Y43_SLICE_X43Y43_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hcccccccc00000000)
  ) CLBLM_R_X27Y43_SLICE_X43Y43_ALUT (
.I0(1'b1),
.I1(CLBLM_R_X27Y43_SLICE_X43Y43_DQ),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLM_R_X27Y43_SLICE_X43Y43_AO5),
.O6(CLBLM_R_X27Y43_SLICE_X43Y43_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT0),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT1),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT2),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT3),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT4),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT5),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X43Y25_IOB_X1Y26_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_BUFGCTRL (
.CE0(CLBLL_L_X24Y46_SLICE_X36Y46_DQ),
.CE1(1'b1),
.I0(RIOB33_X43Y25_IOB_X1Y26_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_O),
.O(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_O),
.O(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_O),
.O(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O),
.O(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y11_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_O),
.O(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y11_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_O),
.O(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y8_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_O),
.O(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y8_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "MMCME2_ADV" *)
  MMCME2_ADV #(
    .BANDWIDTH("OPTIMIZED"),
    .CLKFBOUT_MULT_F(10.750),
    .CLKFBOUT_PHASE(0.000),
    .CLKIN1_PERIOD(11.944),
    .CLKIN2_PERIOD(11.944),
    .CLKOUT0_DIVIDE_F(10.250),
    .CLKOUT0_DUTY_CYCLE(0.500),
    .CLKOUT0_PHASE(43.902),
    .CLKOUT1_DIVIDE(32),
    .CLKOUT1_DUTY_CYCLE(0.5312),
    .CLKOUT1_PHASE(90.000),
    .CLKOUT2_DIVIDE(48),
    .CLKOUT2_DUTY_CYCLE(0.5000),
    .CLKOUT2_PHASE(135.000),
    .CLKOUT3_DIVIDE(64),
    .CLKOUT3_DUTY_CYCLE(0.5000),
    .CLKOUT3_PHASE(45.000),
    .CLKOUT4_DIVIDE(80),
    .CLKOUT4_DUTY_CYCLE(0.5000),
    .CLKOUT4_PHASE(90.000),
    .CLKOUT5_DIVIDE(96),
    .CLKOUT5_DUTY_CYCLE(0.5000),
    .CLKOUT5_PHASE(135.000),
    .CLKOUT6_DIVIDE(1),
    .CLKOUT6_DUTY_CYCLE(0.500),
    .CLKOUT6_PHASE(0.000),
    .COMPENSATION(""),
    .DIVCLK_DIVIDE(1),
    .IS_CLKINSEL_INVERTED(1'b0),
    .IS_PSEN_INVERTED(1'b1),
    .IS_PSINCDEC_INVERTED(1'b1),
    .IS_PWRDWN_INVERTED(1'b0),
    .IS_RST_INVERTED(1'b0),
    .STARTUP_WAIT("FALSE")
  ) CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_MMCME2_ADV (
.CLKFBIN(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBOUT),
.CLKFBOUT(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBOUT),
.CLKFBOUTB(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBOUTB),
.CLKFBSTOPPED(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBSTOPPED),
.CLKIN1(CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y8_O),
.CLKIN2(RIOB33_X43Y25_IOB_X1Y26_I),
.CLKINSEL(LIOB33_X0Y9_IOB_X0Y10_I),
.CLKINSTOPPED(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKINSTOPPED),
.CLKOUT0(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT0),
.CLKOUT0B(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT0B),
.CLKOUT1(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT1),
.CLKOUT1B(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT1B),
.CLKOUT2(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT2),
.CLKOUT2B(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT2B),
.CLKOUT3(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT3),
.CLKOUT3B(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT3B),
.CLKOUT4(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT4),
.CLKOUT5(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT5),
.DADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.DCLK(1'b0),
.DEN(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.DO({CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO15, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO14, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO13, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO12, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO11, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO10, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO9, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO8, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO7, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO6, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO5, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO4, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO3, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO2, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO1, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO0}),
.DRDY(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DRDY),
.DWE(1'b0),
.LOCKED(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_LOCKED),
.PSCLK(1'b0),
.PSDONE(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSDONE),
.PSEN(1'b1),
.PSINCDEC(1'b1),
.PWRDWN(LIOB33_X0Y11_IOB_X0Y12_I),
.RST(CLBLM_R_X27Y8_SLICE_X42Y8_DQ)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y1_OBUF (
.I(LIOB33_X0Y5_IOB_X0Y6_I),
.O(led[7])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y3_IOB_X0Y3_OBUF (
.I(CLBLM_R_X3Y10_SLICE_X2Y10_CQ),
.O(led[0])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y3_IOB_X0Y4_OBUF (
.I(CLBLM_R_X11Y10_SLICE_X15Y10_AQ),
.O(led[5])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y5_IOB_X0Y6_IBUF (
.I(sw[7]),
.O(LIOB33_X0Y5_IOB_X0Y6_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y9_IOB_X0Y10_IBUF (
.I(sw[2]),
.O(LIOB33_X0Y9_IOB_X0Y10_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y11_IOB_X0Y11_IBUF (
.I(sw[0]),
.O(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y11_IOB_X0Y12_IBUF (
.I(sw[1]),
.O(LIOB33_X0Y11_IOB_X0Y12_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y17_IOB_X0Y18_OBUF (
.I(CLBLM_R_X5Y20_SLICE_X7Y20_AQ),
.O(led[4])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y19_IOB_X0Y19_OBUF (
.I(CLBLM_R_X27Y19_SLICE_X43Y19_AQ),
.O(led[3])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y19_IOB_X0Y20_OBUF (
.I(CLBLM_R_X11Y33_SLICE_X14Y33_AQ),
.O(led[2])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y25_IOB_X0Y26_IBUF (
.I(jc4),
.O(LIOB33_X0Y25_IOB_X0Y26_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y27_IOB_X0Y28_OBUF (
.I(LIOB33_X0Y25_IOB_X0Y26_I),
.O(jc2)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y43_IOB_X0Y43_OBUF (
.I(CLBLM_R_X27Y43_SLICE_X43Y43_CQ),
.O(led[1])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y0_IOB_X0Y0_OBUF (
.I(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_LOCKED),
.O(led[6])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y25_IOB_X1Y26_IBUF (
.I(clk),
.O(RIOB33_X43Y25_IOB_X1Y26_I)
  );
  assign CLBLL_L_X24Y46_SLICE_X36Y46_A = CLBLL_L_X24Y46_SLICE_X36Y46_AO6;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_B = CLBLL_L_X24Y46_SLICE_X36Y46_BO6;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_C = CLBLL_L_X24Y46_SLICE_X36Y46_CO6;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_D = CLBLL_L_X24Y46_SLICE_X36Y46_DO6;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_AMUX = CLBLL_L_X24Y46_SLICE_X36Y46_AO6;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_A = CLBLL_L_X24Y46_SLICE_X37Y46_AO6;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_B = CLBLL_L_X24Y46_SLICE_X37Y46_BO6;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_C = CLBLL_L_X24Y46_SLICE_X37Y46_CO6;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_D = CLBLL_L_X24Y46_SLICE_X37Y46_DO6;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_A = CLBLL_L_X26Y9_SLICE_X40Y9_AO6;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_B = CLBLL_L_X26Y9_SLICE_X40Y9_BO6;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_C = CLBLL_L_X26Y9_SLICE_X40Y9_CO6;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_D = CLBLL_L_X26Y9_SLICE_X40Y9_DO6;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_A = CLBLL_L_X26Y9_SLICE_X41Y9_AO6;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_B = CLBLL_L_X26Y9_SLICE_X41Y9_BO6;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_C = CLBLL_L_X26Y9_SLICE_X41Y9_CO6;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_D = CLBLL_L_X26Y9_SLICE_X41Y9_DO6;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_A = CLBLM_R_X3Y5_SLICE_X2Y5_AO6;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_B = CLBLM_R_X3Y5_SLICE_X2Y5_BO6;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_C = CLBLM_R_X3Y5_SLICE_X2Y5_CO6;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_D = CLBLM_R_X3Y5_SLICE_X2Y5_DO6;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_AMUX = CLBLM_R_X3Y5_SLICE_X2Y5_AO6;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_BMUX = CLBLM_R_X3Y5_SLICE_X2Y5_B_XOR;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_CMUX = CLBLM_R_X3Y5_SLICE_X2Y5_C_XOR;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_DMUX = CLBLM_R_X3Y5_SLICE_X2Y5_D_XOR;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_A = CLBLM_R_X3Y5_SLICE_X3Y5_AO6;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_B = CLBLM_R_X3Y5_SLICE_X3Y5_BO6;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_C = CLBLM_R_X3Y5_SLICE_X3Y5_CO6;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_D = CLBLM_R_X3Y5_SLICE_X3Y5_DO6;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_A = CLBLM_R_X3Y6_SLICE_X2Y6_AO6;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_B = CLBLM_R_X3Y6_SLICE_X2Y6_BO6;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_C = CLBLM_R_X3Y6_SLICE_X2Y6_CO6;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_D = CLBLM_R_X3Y6_SLICE_X2Y6_DO6;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_AMUX = CLBLM_R_X3Y6_SLICE_X2Y6_A_XOR;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_BMUX = CLBLM_R_X3Y6_SLICE_X2Y6_B_XOR;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_CMUX = CLBLM_R_X3Y6_SLICE_X2Y6_C_XOR;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_DMUX = CLBLM_R_X3Y6_SLICE_X2Y6_D_XOR;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_A = CLBLM_R_X3Y6_SLICE_X3Y6_AO6;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_B = CLBLM_R_X3Y6_SLICE_X3Y6_BO6;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_C = CLBLM_R_X3Y6_SLICE_X3Y6_CO6;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_D = CLBLM_R_X3Y6_SLICE_X3Y6_DO6;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_A = CLBLM_R_X3Y7_SLICE_X2Y7_AO6;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_B = CLBLM_R_X3Y7_SLICE_X2Y7_BO6;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_C = CLBLM_R_X3Y7_SLICE_X2Y7_CO6;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_D = CLBLM_R_X3Y7_SLICE_X2Y7_DO6;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_AMUX = CLBLM_R_X3Y7_SLICE_X2Y7_A_XOR;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_BMUX = CLBLM_R_X3Y7_SLICE_X2Y7_B_XOR;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_CMUX = CLBLM_R_X3Y7_SLICE_X2Y7_C_XOR;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_DMUX = CLBLM_R_X3Y7_SLICE_X2Y7_D_XOR;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_A = CLBLM_R_X3Y7_SLICE_X3Y7_AO6;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_B = CLBLM_R_X3Y7_SLICE_X3Y7_BO6;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_C = CLBLM_R_X3Y7_SLICE_X3Y7_CO6;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_D = CLBLM_R_X3Y7_SLICE_X3Y7_DO6;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_A = CLBLM_R_X3Y8_SLICE_X2Y8_AO6;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_B = CLBLM_R_X3Y8_SLICE_X2Y8_BO6;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_C = CLBLM_R_X3Y8_SLICE_X2Y8_CO6;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_D = CLBLM_R_X3Y8_SLICE_X2Y8_DO6;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_AMUX = CLBLM_R_X3Y8_SLICE_X2Y8_A5Q;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_BMUX = CLBLM_R_X3Y8_SLICE_X2Y8_B_XOR;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_CMUX = CLBLM_R_X3Y8_SLICE_X2Y8_C_XOR;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_DMUX = CLBLM_R_X3Y8_SLICE_X2Y8_D_XOR;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_A = CLBLM_R_X3Y8_SLICE_X3Y8_AO6;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_B = CLBLM_R_X3Y8_SLICE_X3Y8_BO6;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_C = CLBLM_R_X3Y8_SLICE_X3Y8_CO6;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_D = CLBLM_R_X3Y8_SLICE_X3Y8_DO6;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_A = CLBLM_R_X3Y9_SLICE_X2Y9_AO6;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_B = CLBLM_R_X3Y9_SLICE_X2Y9_BO6;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_C = CLBLM_R_X3Y9_SLICE_X2Y9_CO6;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_D = CLBLM_R_X3Y9_SLICE_X2Y9_DO6;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_AMUX = CLBLM_R_X3Y9_SLICE_X2Y9_A_XOR;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_BMUX = CLBLM_R_X3Y9_SLICE_X2Y9_B_XOR;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_CMUX = CLBLM_R_X3Y9_SLICE_X2Y9_C5Q;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_DMUX = CLBLM_R_X3Y9_SLICE_X2Y9_D_XOR;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_A = CLBLM_R_X3Y9_SLICE_X3Y9_AO6;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_B = CLBLM_R_X3Y9_SLICE_X3Y9_BO6;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_C = CLBLM_R_X3Y9_SLICE_X3Y9_CO6;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_D = CLBLM_R_X3Y9_SLICE_X3Y9_DO6;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_A = CLBLM_R_X3Y10_SLICE_X2Y10_AO6;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_B = CLBLM_R_X3Y10_SLICE_X2Y10_BO6;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_C = CLBLM_R_X3Y10_SLICE_X2Y10_CO6;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_D = CLBLM_R_X3Y10_SLICE_X2Y10_DO6;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_AMUX = CLBLM_R_X3Y10_SLICE_X2Y10_A_XOR;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_BMUX = CLBLM_R_X3Y10_SLICE_X2Y10_B_XOR;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_CMUX = CLBLM_R_X3Y10_SLICE_X2Y10_C_XOR;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_DMUX = CLBLM_R_X3Y10_SLICE_X2Y10_D_XOR;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_A = CLBLM_R_X3Y10_SLICE_X3Y10_AO6;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_B = CLBLM_R_X3Y10_SLICE_X3Y10_BO6;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_C = CLBLM_R_X3Y10_SLICE_X3Y10_CO6;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_D = CLBLM_R_X3Y10_SLICE_X3Y10_DO6;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_A = CLBLM_R_X5Y15_SLICE_X6Y15_AO6;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_B = CLBLM_R_X5Y15_SLICE_X6Y15_BO6;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_C = CLBLM_R_X5Y15_SLICE_X6Y15_CO6;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_D = CLBLM_R_X5Y15_SLICE_X6Y15_DO6;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_A = CLBLM_R_X5Y15_SLICE_X7Y15_AO6;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_B = CLBLM_R_X5Y15_SLICE_X7Y15_BO6;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_C = CLBLM_R_X5Y15_SLICE_X7Y15_CO6;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_D = CLBLM_R_X5Y15_SLICE_X7Y15_DO6;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_AMUX = CLBLM_R_X5Y15_SLICE_X7Y15_AO6;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_BMUX = CLBLM_R_X5Y15_SLICE_X7Y15_B_XOR;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_CMUX = CLBLM_R_X5Y15_SLICE_X7Y15_C_XOR;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_DMUX = CLBLM_R_X5Y15_SLICE_X7Y15_D_XOR;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_A = CLBLM_R_X5Y16_SLICE_X6Y16_AO6;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_B = CLBLM_R_X5Y16_SLICE_X6Y16_BO6;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_C = CLBLM_R_X5Y16_SLICE_X6Y16_CO6;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_D = CLBLM_R_X5Y16_SLICE_X6Y16_DO6;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_A = CLBLM_R_X5Y16_SLICE_X7Y16_AO6;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_B = CLBLM_R_X5Y16_SLICE_X7Y16_BO6;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_C = CLBLM_R_X5Y16_SLICE_X7Y16_CO6;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_D = CLBLM_R_X5Y16_SLICE_X7Y16_DO6;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_AMUX = CLBLM_R_X5Y16_SLICE_X7Y16_A_XOR;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_BMUX = CLBLM_R_X5Y16_SLICE_X7Y16_B_XOR;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_CMUX = CLBLM_R_X5Y16_SLICE_X7Y16_C_XOR;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_DMUX = CLBLM_R_X5Y16_SLICE_X7Y16_D_XOR;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_A = CLBLM_R_X5Y17_SLICE_X6Y17_AO6;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_B = CLBLM_R_X5Y17_SLICE_X6Y17_BO6;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_C = CLBLM_R_X5Y17_SLICE_X6Y17_CO6;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_D = CLBLM_R_X5Y17_SLICE_X6Y17_DO6;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_A = CLBLM_R_X5Y17_SLICE_X7Y17_AO6;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_B = CLBLM_R_X5Y17_SLICE_X7Y17_BO6;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_C = CLBLM_R_X5Y17_SLICE_X7Y17_CO6;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_D = CLBLM_R_X5Y17_SLICE_X7Y17_DO6;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_AMUX = CLBLM_R_X5Y17_SLICE_X7Y17_A_XOR;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_BMUX = CLBLM_R_X5Y17_SLICE_X7Y17_B_XOR;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_CMUX = CLBLM_R_X5Y17_SLICE_X7Y17_C_XOR;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_DMUX = CLBLM_R_X5Y17_SLICE_X7Y17_D_XOR;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_A = CLBLM_R_X5Y18_SLICE_X6Y18_AO6;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_B = CLBLM_R_X5Y18_SLICE_X6Y18_BO6;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_C = CLBLM_R_X5Y18_SLICE_X6Y18_CO6;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_D = CLBLM_R_X5Y18_SLICE_X6Y18_DO6;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_A = CLBLM_R_X5Y18_SLICE_X7Y18_AO6;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_B = CLBLM_R_X5Y18_SLICE_X7Y18_BO6;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_C = CLBLM_R_X5Y18_SLICE_X7Y18_CO6;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_D = CLBLM_R_X5Y18_SLICE_X7Y18_DO6;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_BMUX = CLBLM_R_X5Y18_SLICE_X7Y18_B_XOR;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_CMUX = CLBLM_R_X5Y18_SLICE_X7Y18_C_XOR;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_DMUX = CLBLM_R_X5Y18_SLICE_X7Y18_D_XOR;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_A = CLBLM_R_X5Y19_SLICE_X6Y19_AO6;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_B = CLBLM_R_X5Y19_SLICE_X6Y19_BO6;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_C = CLBLM_R_X5Y19_SLICE_X6Y19_CO6;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_D = CLBLM_R_X5Y19_SLICE_X6Y19_DO6;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_A = CLBLM_R_X5Y19_SLICE_X7Y19_AO6;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_B = CLBLM_R_X5Y19_SLICE_X7Y19_BO6;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_C = CLBLM_R_X5Y19_SLICE_X7Y19_CO6;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_D = CLBLM_R_X5Y19_SLICE_X7Y19_DO6;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_BMUX = CLBLM_R_X5Y19_SLICE_X7Y19_B_XOR;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_CMUX = CLBLM_R_X5Y19_SLICE_X7Y19_C_XOR;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_DMUX = CLBLM_R_X5Y19_SLICE_X7Y19_D_XOR;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_A = CLBLM_R_X5Y20_SLICE_X6Y20_AO6;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_B = CLBLM_R_X5Y20_SLICE_X6Y20_BO6;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_C = CLBLM_R_X5Y20_SLICE_X6Y20_CO6;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_D = CLBLM_R_X5Y20_SLICE_X6Y20_DO6;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_A = CLBLM_R_X5Y20_SLICE_X7Y20_AO6;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_B = CLBLM_R_X5Y20_SLICE_X7Y20_BO6;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_C = CLBLM_R_X5Y20_SLICE_X7Y20_CO6;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_D = CLBLM_R_X5Y20_SLICE_X7Y20_DO6;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_AMUX = CLBLM_R_X5Y20_SLICE_X7Y20_A_XOR;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_BMUX = CLBLM_R_X5Y20_SLICE_X7Y20_B_XOR;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_A = CLBLM_R_X11Y5_SLICE_X14Y5_AO6;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_B = CLBLM_R_X11Y5_SLICE_X14Y5_BO6;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_C = CLBLM_R_X11Y5_SLICE_X14Y5_CO6;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_D = CLBLM_R_X11Y5_SLICE_X14Y5_DO6;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_A = CLBLM_R_X11Y5_SLICE_X15Y5_AO6;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_B = CLBLM_R_X11Y5_SLICE_X15Y5_BO6;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_C = CLBLM_R_X11Y5_SLICE_X15Y5_CO6;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_D = CLBLM_R_X11Y5_SLICE_X15Y5_DO6;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_AMUX = CLBLM_R_X11Y5_SLICE_X15Y5_AO6;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_BMUX = CLBLM_R_X11Y5_SLICE_X15Y5_B_XOR;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_CMUX = CLBLM_R_X11Y5_SLICE_X15Y5_C_XOR;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_DMUX = CLBLM_R_X11Y5_SLICE_X15Y5_D_XOR;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_A = CLBLM_R_X11Y6_SLICE_X14Y6_AO6;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_B = CLBLM_R_X11Y6_SLICE_X14Y6_BO6;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_C = CLBLM_R_X11Y6_SLICE_X14Y6_CO6;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_D = CLBLM_R_X11Y6_SLICE_X14Y6_DO6;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_A = CLBLM_R_X11Y6_SLICE_X15Y6_AO6;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_B = CLBLM_R_X11Y6_SLICE_X15Y6_BO6;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_C = CLBLM_R_X11Y6_SLICE_X15Y6_CO6;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_D = CLBLM_R_X11Y6_SLICE_X15Y6_DO6;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_AMUX = CLBLM_R_X11Y6_SLICE_X15Y6_A_XOR;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_BMUX = CLBLM_R_X11Y6_SLICE_X15Y6_B_XOR;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_CMUX = CLBLM_R_X11Y6_SLICE_X15Y6_C_XOR;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_DMUX = CLBLM_R_X11Y6_SLICE_X15Y6_D_XOR;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_A = CLBLM_R_X11Y7_SLICE_X14Y7_AO6;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_B = CLBLM_R_X11Y7_SLICE_X14Y7_BO6;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_C = CLBLM_R_X11Y7_SLICE_X14Y7_CO6;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_D = CLBLM_R_X11Y7_SLICE_X14Y7_DO6;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_A = CLBLM_R_X11Y7_SLICE_X15Y7_AO6;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_B = CLBLM_R_X11Y7_SLICE_X15Y7_BO6;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_C = CLBLM_R_X11Y7_SLICE_X15Y7_CO6;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_D = CLBLM_R_X11Y7_SLICE_X15Y7_DO6;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_AMUX = CLBLM_R_X11Y7_SLICE_X15Y7_A_XOR;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_BMUX = CLBLM_R_X11Y7_SLICE_X15Y7_B_XOR;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_CMUX = CLBLM_R_X11Y7_SLICE_X15Y7_C_XOR;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_DMUX = CLBLM_R_X11Y7_SLICE_X15Y7_D_XOR;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_A = CLBLM_R_X11Y8_SLICE_X14Y8_AO6;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_B = CLBLM_R_X11Y8_SLICE_X14Y8_BO6;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_C = CLBLM_R_X11Y8_SLICE_X14Y8_CO6;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_D = CLBLM_R_X11Y8_SLICE_X14Y8_DO6;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_A = CLBLM_R_X11Y8_SLICE_X15Y8_AO6;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_B = CLBLM_R_X11Y8_SLICE_X15Y8_BO6;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_C = CLBLM_R_X11Y8_SLICE_X15Y8_CO6;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_D = CLBLM_R_X11Y8_SLICE_X15Y8_DO6;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_BMUX = CLBLM_R_X11Y8_SLICE_X15Y8_B_XOR;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_CMUX = CLBLM_R_X11Y8_SLICE_X15Y8_C_XOR;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_DMUX = CLBLM_R_X11Y8_SLICE_X15Y8_D_XOR;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_A = CLBLM_R_X11Y9_SLICE_X14Y9_AO6;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_B = CLBLM_R_X11Y9_SLICE_X14Y9_BO6;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_C = CLBLM_R_X11Y9_SLICE_X14Y9_CO6;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_D = CLBLM_R_X11Y9_SLICE_X14Y9_DO6;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_A = CLBLM_R_X11Y9_SLICE_X15Y9_AO6;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_B = CLBLM_R_X11Y9_SLICE_X15Y9_BO6;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_C = CLBLM_R_X11Y9_SLICE_X15Y9_CO6;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_D = CLBLM_R_X11Y9_SLICE_X15Y9_DO6;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_BMUX = CLBLM_R_X11Y9_SLICE_X15Y9_B_XOR;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_CMUX = CLBLM_R_X11Y9_SLICE_X15Y9_C_XOR;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_DMUX = CLBLM_R_X11Y9_SLICE_X15Y9_D_XOR;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_A = CLBLM_R_X11Y10_SLICE_X14Y10_AO6;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_B = CLBLM_R_X11Y10_SLICE_X14Y10_BO6;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_C = CLBLM_R_X11Y10_SLICE_X14Y10_CO6;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_D = CLBLM_R_X11Y10_SLICE_X14Y10_DO6;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_A = CLBLM_R_X11Y10_SLICE_X15Y10_AO6;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_B = CLBLM_R_X11Y10_SLICE_X15Y10_BO6;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_C = CLBLM_R_X11Y10_SLICE_X15Y10_CO6;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_D = CLBLM_R_X11Y10_SLICE_X15Y10_DO6;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_AMUX = CLBLM_R_X11Y10_SLICE_X15Y10_A_XOR;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_BMUX = CLBLM_R_X11Y10_SLICE_X15Y10_B_XOR;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_A = CLBLM_R_X11Y28_SLICE_X14Y28_AO6;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_B = CLBLM_R_X11Y28_SLICE_X14Y28_BO6;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_C = CLBLM_R_X11Y28_SLICE_X14Y28_CO6;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_D = CLBLM_R_X11Y28_SLICE_X14Y28_DO6;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_AMUX = CLBLM_R_X11Y28_SLICE_X14Y28_AO6;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_BMUX = CLBLM_R_X11Y28_SLICE_X14Y28_B_XOR;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_CMUX = CLBLM_R_X11Y28_SLICE_X14Y28_C_XOR;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_DMUX = CLBLM_R_X11Y28_SLICE_X14Y28_D_XOR;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_A = CLBLM_R_X11Y28_SLICE_X15Y28_AO6;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_B = CLBLM_R_X11Y28_SLICE_X15Y28_BO6;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_C = CLBLM_R_X11Y28_SLICE_X15Y28_CO6;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_D = CLBLM_R_X11Y28_SLICE_X15Y28_DO6;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_A = CLBLM_R_X11Y29_SLICE_X14Y29_AO6;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_B = CLBLM_R_X11Y29_SLICE_X14Y29_BO6;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_C = CLBLM_R_X11Y29_SLICE_X14Y29_CO6;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_D = CLBLM_R_X11Y29_SLICE_X14Y29_DO6;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_AMUX = CLBLM_R_X11Y29_SLICE_X14Y29_A_XOR;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_BMUX = CLBLM_R_X11Y29_SLICE_X14Y29_B_XOR;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_CMUX = CLBLM_R_X11Y29_SLICE_X14Y29_C_XOR;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_DMUX = CLBLM_R_X11Y29_SLICE_X14Y29_D_XOR;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_A = CLBLM_R_X11Y29_SLICE_X15Y29_AO6;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_B = CLBLM_R_X11Y29_SLICE_X15Y29_BO6;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_C = CLBLM_R_X11Y29_SLICE_X15Y29_CO6;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_D = CLBLM_R_X11Y29_SLICE_X15Y29_DO6;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_A = CLBLM_R_X11Y30_SLICE_X14Y30_AO6;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_B = CLBLM_R_X11Y30_SLICE_X14Y30_BO6;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_C = CLBLM_R_X11Y30_SLICE_X14Y30_CO6;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_D = CLBLM_R_X11Y30_SLICE_X14Y30_DO6;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_AMUX = CLBLM_R_X11Y30_SLICE_X14Y30_A_XOR;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_BMUX = CLBLM_R_X11Y30_SLICE_X14Y30_B_XOR;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_CMUX = CLBLM_R_X11Y30_SLICE_X14Y30_C_XOR;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_DMUX = CLBLM_R_X11Y30_SLICE_X14Y30_D_XOR;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_A = CLBLM_R_X11Y30_SLICE_X15Y30_AO6;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_B = CLBLM_R_X11Y30_SLICE_X15Y30_BO6;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_C = CLBLM_R_X11Y30_SLICE_X15Y30_CO6;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_D = CLBLM_R_X11Y30_SLICE_X15Y30_DO6;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_A = CLBLM_R_X11Y31_SLICE_X14Y31_AO6;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_B = CLBLM_R_X11Y31_SLICE_X14Y31_BO6;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_C = CLBLM_R_X11Y31_SLICE_X14Y31_CO6;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_D = CLBLM_R_X11Y31_SLICE_X14Y31_DO6;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_BMUX = CLBLM_R_X11Y31_SLICE_X14Y31_B_XOR;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_CMUX = CLBLM_R_X11Y31_SLICE_X14Y31_C_XOR;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_DMUX = CLBLM_R_X11Y31_SLICE_X14Y31_D_XOR;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_A = CLBLM_R_X11Y31_SLICE_X15Y31_AO6;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_B = CLBLM_R_X11Y31_SLICE_X15Y31_BO6;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_C = CLBLM_R_X11Y31_SLICE_X15Y31_CO6;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_D = CLBLM_R_X11Y31_SLICE_X15Y31_DO6;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_A = CLBLM_R_X11Y32_SLICE_X14Y32_AO6;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_B = CLBLM_R_X11Y32_SLICE_X14Y32_BO6;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_C = CLBLM_R_X11Y32_SLICE_X14Y32_CO6;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_D = CLBLM_R_X11Y32_SLICE_X14Y32_DO6;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_BMUX = CLBLM_R_X11Y32_SLICE_X14Y32_B_XOR;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_CMUX = CLBLM_R_X11Y32_SLICE_X14Y32_C_XOR;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_DMUX = CLBLM_R_X11Y32_SLICE_X14Y32_D_XOR;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_A = CLBLM_R_X11Y32_SLICE_X15Y32_AO6;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_B = CLBLM_R_X11Y32_SLICE_X15Y32_BO6;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_C = CLBLM_R_X11Y32_SLICE_X15Y32_CO6;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_D = CLBLM_R_X11Y32_SLICE_X15Y32_DO6;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_A = CLBLM_R_X11Y33_SLICE_X14Y33_AO6;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_B = CLBLM_R_X11Y33_SLICE_X14Y33_BO6;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_C = CLBLM_R_X11Y33_SLICE_X14Y33_CO6;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_D = CLBLM_R_X11Y33_SLICE_X14Y33_DO6;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_AMUX = CLBLM_R_X11Y33_SLICE_X14Y33_A_XOR;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_BMUX = CLBLM_R_X11Y33_SLICE_X14Y33_B_XOR;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_A = CLBLM_R_X11Y33_SLICE_X15Y33_AO6;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_B = CLBLM_R_X11Y33_SLICE_X15Y33_BO6;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_C = CLBLM_R_X11Y33_SLICE_X15Y33_CO6;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_D = CLBLM_R_X11Y33_SLICE_X15Y33_DO6;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_A = CLBLM_R_X27Y8_SLICE_X42Y8_AO6;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_B = CLBLM_R_X27Y8_SLICE_X42Y8_BO6;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_C = CLBLM_R_X27Y8_SLICE_X42Y8_CO6;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_D = CLBLM_R_X27Y8_SLICE_X42Y8_DO6;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_A = CLBLM_R_X27Y8_SLICE_X43Y8_AO6;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_B = CLBLM_R_X27Y8_SLICE_X43Y8_BO6;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_C = CLBLM_R_X27Y8_SLICE_X43Y8_CO6;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_D = CLBLM_R_X27Y8_SLICE_X43Y8_DO6;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_A = CLBLM_R_X27Y14_SLICE_X42Y14_AO6;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_B = CLBLM_R_X27Y14_SLICE_X42Y14_BO6;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_C = CLBLM_R_X27Y14_SLICE_X42Y14_CO6;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_D = CLBLM_R_X27Y14_SLICE_X42Y14_DO6;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_A = CLBLM_R_X27Y14_SLICE_X43Y14_AO6;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_B = CLBLM_R_X27Y14_SLICE_X43Y14_BO6;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_C = CLBLM_R_X27Y14_SLICE_X43Y14_CO6;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_D = CLBLM_R_X27Y14_SLICE_X43Y14_DO6;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_AMUX = CLBLM_R_X27Y14_SLICE_X43Y14_AO6;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_BMUX = CLBLM_R_X27Y14_SLICE_X43Y14_B_XOR;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_CMUX = CLBLM_R_X27Y14_SLICE_X43Y14_C_XOR;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_DMUX = CLBLM_R_X27Y14_SLICE_X43Y14_D_XOR;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_A = CLBLM_R_X27Y15_SLICE_X42Y15_AO6;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_B = CLBLM_R_X27Y15_SLICE_X42Y15_BO6;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_C = CLBLM_R_X27Y15_SLICE_X42Y15_CO6;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_D = CLBLM_R_X27Y15_SLICE_X42Y15_DO6;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_A = CLBLM_R_X27Y15_SLICE_X43Y15_AO6;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_B = CLBLM_R_X27Y15_SLICE_X43Y15_BO6;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_C = CLBLM_R_X27Y15_SLICE_X43Y15_CO6;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_D = CLBLM_R_X27Y15_SLICE_X43Y15_DO6;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_AMUX = CLBLM_R_X27Y15_SLICE_X43Y15_A_XOR;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_BMUX = CLBLM_R_X27Y15_SLICE_X43Y15_B_XOR;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_CMUX = CLBLM_R_X27Y15_SLICE_X43Y15_C_XOR;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_DMUX = CLBLM_R_X27Y15_SLICE_X43Y15_D_XOR;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_A = CLBLM_R_X27Y16_SLICE_X42Y16_AO6;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_B = CLBLM_R_X27Y16_SLICE_X42Y16_BO6;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_C = CLBLM_R_X27Y16_SLICE_X42Y16_CO6;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_D = CLBLM_R_X27Y16_SLICE_X42Y16_DO6;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_A = CLBLM_R_X27Y16_SLICE_X43Y16_AO6;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_B = CLBLM_R_X27Y16_SLICE_X43Y16_BO6;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_C = CLBLM_R_X27Y16_SLICE_X43Y16_CO6;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_D = CLBLM_R_X27Y16_SLICE_X43Y16_DO6;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_AMUX = CLBLM_R_X27Y16_SLICE_X43Y16_A_XOR;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_BMUX = CLBLM_R_X27Y16_SLICE_X43Y16_B_XOR;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_CMUX = CLBLM_R_X27Y16_SLICE_X43Y16_C_XOR;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_DMUX = CLBLM_R_X27Y16_SLICE_X43Y16_D_XOR;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_A = CLBLM_R_X27Y17_SLICE_X42Y17_AO6;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_B = CLBLM_R_X27Y17_SLICE_X42Y17_BO6;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_C = CLBLM_R_X27Y17_SLICE_X42Y17_CO6;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_D = CLBLM_R_X27Y17_SLICE_X42Y17_DO6;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_A = CLBLM_R_X27Y17_SLICE_X43Y17_AO6;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_B = CLBLM_R_X27Y17_SLICE_X43Y17_BO6;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_C = CLBLM_R_X27Y17_SLICE_X43Y17_CO6;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_D = CLBLM_R_X27Y17_SLICE_X43Y17_DO6;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_BMUX = CLBLM_R_X27Y17_SLICE_X43Y17_B_XOR;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_CMUX = CLBLM_R_X27Y17_SLICE_X43Y17_C_XOR;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_DMUX = CLBLM_R_X27Y17_SLICE_X43Y17_D_XOR;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_A = CLBLM_R_X27Y18_SLICE_X42Y18_AO6;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_B = CLBLM_R_X27Y18_SLICE_X42Y18_BO6;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_C = CLBLM_R_X27Y18_SLICE_X42Y18_CO6;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_D = CLBLM_R_X27Y18_SLICE_X42Y18_DO6;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_A = CLBLM_R_X27Y18_SLICE_X43Y18_AO6;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_B = CLBLM_R_X27Y18_SLICE_X43Y18_BO6;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_C = CLBLM_R_X27Y18_SLICE_X43Y18_CO6;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_D = CLBLM_R_X27Y18_SLICE_X43Y18_DO6;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_BMUX = CLBLM_R_X27Y18_SLICE_X43Y18_B_XOR;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_CMUX = CLBLM_R_X27Y18_SLICE_X43Y18_C_XOR;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_DMUX = CLBLM_R_X27Y18_SLICE_X43Y18_D_XOR;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_A = CLBLM_R_X27Y19_SLICE_X42Y19_AO6;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_B = CLBLM_R_X27Y19_SLICE_X42Y19_BO6;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_C = CLBLM_R_X27Y19_SLICE_X42Y19_CO6;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_D = CLBLM_R_X27Y19_SLICE_X42Y19_DO6;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_A = CLBLM_R_X27Y19_SLICE_X43Y19_AO6;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_B = CLBLM_R_X27Y19_SLICE_X43Y19_BO6;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_C = CLBLM_R_X27Y19_SLICE_X43Y19_CO6;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_D = CLBLM_R_X27Y19_SLICE_X43Y19_DO6;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_AMUX = CLBLM_R_X27Y19_SLICE_X43Y19_A_XOR;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_BMUX = CLBLM_R_X27Y19_SLICE_X43Y19_B_XOR;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_CMUX = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_A = CLBLM_R_X27Y38_SLICE_X42Y38_AO6;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_B = CLBLM_R_X27Y38_SLICE_X42Y38_BO6;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_C = CLBLM_R_X27Y38_SLICE_X42Y38_CO6;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_D = CLBLM_R_X27Y38_SLICE_X42Y38_DO6;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_A = CLBLM_R_X27Y38_SLICE_X43Y38_AO6;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_B = CLBLM_R_X27Y38_SLICE_X43Y38_BO6;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_C = CLBLM_R_X27Y38_SLICE_X43Y38_CO6;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_D = CLBLM_R_X27Y38_SLICE_X43Y38_DO6;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_AMUX = CLBLM_R_X27Y38_SLICE_X43Y38_AO6;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_BMUX = CLBLM_R_X27Y38_SLICE_X43Y38_B_XOR;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_CMUX = CLBLM_R_X27Y38_SLICE_X43Y38_C_XOR;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_DMUX = CLBLM_R_X27Y38_SLICE_X43Y38_D_XOR;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_A = CLBLM_R_X27Y39_SLICE_X42Y39_AO6;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_B = CLBLM_R_X27Y39_SLICE_X42Y39_BO6;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_C = CLBLM_R_X27Y39_SLICE_X42Y39_CO6;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_D = CLBLM_R_X27Y39_SLICE_X42Y39_DO6;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_A = CLBLM_R_X27Y39_SLICE_X43Y39_AO6;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_B = CLBLM_R_X27Y39_SLICE_X43Y39_BO6;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_C = CLBLM_R_X27Y39_SLICE_X43Y39_CO6;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_D = CLBLM_R_X27Y39_SLICE_X43Y39_DO6;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_AMUX = CLBLM_R_X27Y39_SLICE_X43Y39_A_XOR;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_BMUX = CLBLM_R_X27Y39_SLICE_X43Y39_B_XOR;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_CMUX = CLBLM_R_X27Y39_SLICE_X43Y39_C_XOR;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_DMUX = CLBLM_R_X27Y39_SLICE_X43Y39_D_XOR;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_A = CLBLM_R_X27Y40_SLICE_X42Y40_AO6;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_B = CLBLM_R_X27Y40_SLICE_X42Y40_BO6;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_C = CLBLM_R_X27Y40_SLICE_X42Y40_CO6;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_D = CLBLM_R_X27Y40_SLICE_X42Y40_DO6;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_A = CLBLM_R_X27Y40_SLICE_X43Y40_AO6;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_B = CLBLM_R_X27Y40_SLICE_X43Y40_BO6;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_C = CLBLM_R_X27Y40_SLICE_X43Y40_CO6;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_D = CLBLM_R_X27Y40_SLICE_X43Y40_DO6;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_AMUX = CLBLM_R_X27Y40_SLICE_X43Y40_A_XOR;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_BMUX = CLBLM_R_X27Y40_SLICE_X43Y40_B_XOR;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_CMUX = CLBLM_R_X27Y40_SLICE_X43Y40_C_XOR;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_DMUX = CLBLM_R_X27Y40_SLICE_X43Y40_D_XOR;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_A = CLBLM_R_X27Y41_SLICE_X42Y41_AO6;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_B = CLBLM_R_X27Y41_SLICE_X42Y41_BO6;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_C = CLBLM_R_X27Y41_SLICE_X42Y41_CO6;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_D = CLBLM_R_X27Y41_SLICE_X42Y41_DO6;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_A = CLBLM_R_X27Y41_SLICE_X43Y41_AO6;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_B = CLBLM_R_X27Y41_SLICE_X43Y41_BO6;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_C = CLBLM_R_X27Y41_SLICE_X43Y41_CO6;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_D = CLBLM_R_X27Y41_SLICE_X43Y41_DO6;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_AMUX = CLBLM_R_X27Y41_SLICE_X43Y41_A5Q;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_BMUX = CLBLM_R_X27Y41_SLICE_X43Y41_B_XOR;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_CMUX = CLBLM_R_X27Y41_SLICE_X43Y41_C_XOR;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_DMUX = CLBLM_R_X27Y41_SLICE_X43Y41_D_XOR;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_A = CLBLM_R_X27Y42_SLICE_X42Y42_AO6;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_B = CLBLM_R_X27Y42_SLICE_X42Y42_BO6;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_C = CLBLM_R_X27Y42_SLICE_X42Y42_CO6;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_D = CLBLM_R_X27Y42_SLICE_X42Y42_DO6;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_A = CLBLM_R_X27Y42_SLICE_X43Y42_AO6;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_B = CLBLM_R_X27Y42_SLICE_X43Y42_BO6;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_C = CLBLM_R_X27Y42_SLICE_X43Y42_CO6;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_D = CLBLM_R_X27Y42_SLICE_X43Y42_DO6;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_AMUX = CLBLM_R_X27Y42_SLICE_X43Y42_A5Q;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_BMUX = CLBLM_R_X27Y42_SLICE_X43Y42_B_XOR;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_CMUX = CLBLM_R_X27Y42_SLICE_X43Y42_C_XOR;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_DMUX = CLBLM_R_X27Y42_SLICE_X43Y42_D_XOR;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_A = CLBLM_R_X27Y43_SLICE_X42Y43_AO6;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_B = CLBLM_R_X27Y43_SLICE_X42Y43_BO6;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_C = CLBLM_R_X27Y43_SLICE_X42Y43_CO6;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_D = CLBLM_R_X27Y43_SLICE_X42Y43_DO6;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_A = CLBLM_R_X27Y43_SLICE_X43Y43_AO6;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_B = CLBLM_R_X27Y43_SLICE_X43Y43_BO6;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_C = CLBLM_R_X27Y43_SLICE_X43Y43_CO6;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_D = CLBLM_R_X27Y43_SLICE_X43Y43_DO6;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_AMUX = CLBLM_R_X27Y43_SLICE_X43Y43_A_XOR;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_BMUX = CLBLM_R_X27Y43_SLICE_X43Y43_B_XOR;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_CMUX = CLBLM_R_X27Y43_SLICE_X43Y43_C_XOR;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_DMUX = CLBLM_R_X27Y43_SLICE_X43Y43_D_XOR;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_OQ = LIOB33_X0Y5_IOB_X0Y6_I;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_TQ = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_OQ = CLBLM_R_X11Y10_SLICE_X15Y10_AQ;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_TQ = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_OQ = CLBLM_R_X3Y10_SLICE_X2Y10_CQ;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_TQ = 1'b1;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_O = LIOB33_X0Y5_IOB_X0Y6_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_O = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_O = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_O = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_OQ = CLBLM_R_X5Y20_SLICE_X7Y20_AQ;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_TQ = 1'b1;
  assign LIOI3_X0Y25_ILOGIC_X0Y26_O = LIOB33_X0Y25_IOB_X0Y26_I;
  assign LIOI3_X0Y27_OLOGIC_X0Y28_OQ = LIOB33_X0Y25_IOB_X0Y26_I;
  assign LIOI3_X0Y27_OLOGIC_X0Y28_TQ = 1'b1;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_OQ = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_LOCKED;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_OQ = CLBLM_R_X11Y33_SLICE_X14Y33_AQ;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_OQ = CLBLM_R_X27Y19_SLICE_X43Y19_AQ;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ = CLBLM_R_X27Y43_SLICE_X43Y43_CQ;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ = 1'b1;
  assign RIOI3_X43Y25_ILOGIC_X1Y26_O = RIOB33_X43Y25_IOB_X1Y26_I;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_D2 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_B6 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_D3 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_D1 = CLBLM_R_X11Y33_SLICE_X14Y33_AQ;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_D4 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_A3 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_D5 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_D5 = CLBLM_R_X27Y14_SLICE_X43Y14_BQ;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_D6 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_A1 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_A2 = CLBLM_R_X11Y31_SLICE_X14Y31_AQ;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_A3 = 1'b1;
  assign LIOB33_X0Y1_IOB_X0Y1_O = LIOB33_X0Y5_IOB_X0Y6_I;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_A4 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_A5 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_A6 = 1'b1;
  assign LIOI3_X0Y25_ILOGIC_X0Y26_D = LIOB33_X0Y25_IOB_X0Y26_I;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_T1 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_AX = 1'b0;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_B1 = CLBLM_R_X11Y31_SLICE_X14Y31_C_XOR;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_C2 = CLBLM_R_X27Y18_SLICE_X43Y18_D_XOR;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_B2 = CLBLM_R_X11Y31_SLICE_X14Y31_DQ;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_C3 = CLBLM_R_X27Y18_SLICE_X43Y18_BQ;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_B3 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_C4 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_B4 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_C5 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_B5 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_C6 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_B6 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_A1 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_A1 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_A2 = CLBLM_R_X11Y10_SLICE_X15Y10_BQ;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_A3 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_A4 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_A5 = CLBLM_R_X11Y10_SLICE_X15Y10_B_XOR;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_A6 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_CIN = CLBLM_R_X27Y17_SLICE_X43Y17_COUT;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_B1 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_AX = 1'b0;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_B1 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_B2 = CLBLM_R_X11Y10_SLICE_X15Y10_AQ;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_B3 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_B4 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_B5 = CLBLM_R_X11Y10_SLICE_X15Y10_A_XOR;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_B6 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_BX = 1'b0;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_BX = 1'b0;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_D1 = CLBLM_R_X27Y19_SLICE_X43Y19_AQ;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_C1 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_C2 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_C3 = CLBLM_R_X11Y10_SLICE_X15Y10_CQ;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_C4 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_C5 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_C6 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_C1 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_CIN = CLBLM_R_X11Y9_SLICE_X15Y9_COUT;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_A2 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_B2 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_C2 = CLBLM_R_X11Y31_SLICE_X14Y31_D_XOR;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_CX = 1'b0;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_D6 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_A1 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_A2 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_A3 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_A4 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_A5 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_A6 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_D1 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_D2 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_D3 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_B1 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_B2 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_B3 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_B4 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_B5 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_B6 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_A1 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_A2 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_A3 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_C1 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_C2 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_C3 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_C4 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_C5 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_C6 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_A5 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_A6 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_B1 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_B2 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_B3 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_B4 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_B5 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_D1 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_D2 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_D3 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_D4 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_D5 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X3Y5_D6 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_C1 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_C2 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_C3 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_C4 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_C5 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_A1 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_A2 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_A3 = CLBLM_R_X3Y5_SLICE_X2Y5_DQ;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_A4 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_A5 = CLBLM_R_X3Y5_SLICE_X2Y5_C_XOR;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_A6 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_D1 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_D2 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_AX = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_D3 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_B1 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_B2 = CLBLM_R_X3Y5_SLICE_X2Y5_CQ;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_B3 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_B4 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_B5 = CLBLM_R_X3Y5_SLICE_X2Y5_D_XOR;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_B6 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_D6 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_CX = 1'b0;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_BX = 1'b0;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_A5 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_C1 = CLBLM_R_X3Y5_SLICE_X2Y5_AQ;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_C2 = CLBLM_R_X3Y5_SLICE_X2Y5_B_XOR;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_C3 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_C4 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_C5 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_C6 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_D1 = CLBLM_R_X11Y31_SLICE_X14Y31_B_XOR;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_D2 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_B4 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_A1 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_D3 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_A2 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_CX = 1'b0;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_A3 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_D1 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_D2 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_D3 = CLBLM_R_X3Y5_SLICE_X2Y5_AO6;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_D4 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_D5 = CLBLM_R_X3Y5_SLICE_X2Y5_BQ;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_D6 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_D4 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_D5 = CLBLM_R_X11Y31_SLICE_X14Y31_CQ;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_A4 = 1'b1;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_DX = 1'b0;
  assign CLBLM_R_X3Y5_SLICE_X2Y5_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_D6 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_A5 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_A6 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_B5 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_B6 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_B1 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_B2 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_B3 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_B4 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_B5 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_B6 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S1 = 1'b1;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_D = LIOB33_X0Y5_IOB_X0Y6_I;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_B3 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_C1 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_B4 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_C2 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_C3 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_C4 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_C5 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_CE1 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_C6 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_S1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_S1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_S1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_CE0 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_C3 = CLBLM_R_X11Y32_SLICE_X14Y32_BQ;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_A1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_S1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_CE0 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_B1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_S1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_S1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_CE0 = CLBLL_L_X24Y46_SLICE_X36Y46_DQ;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_CE1 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_C1 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_A2 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_CIN = CLBLM_R_X5Y15_SLICE_X7Y15_COUT;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_B2 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_D1 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_D2 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_C2 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_D3 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_A3 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_D4 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_D5 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_B3 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X42Y18_D6 = 1'b1;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_D1 = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_LOCKED;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_C3 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_A4 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_D3 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_B4 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_A1 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_A2 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_A3 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_A4 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_A5 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_A6 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_B1 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_B2 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_B3 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_B4 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_B5 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_B6 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_D6 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_C4 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_A5 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_C1 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_C2 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_C3 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_C4 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_C5 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_C6 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_DX = 1'b0;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_B5 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_D1 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_D2 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_D3 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_D4 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_D5 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X3Y6_D6 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_C4 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_C5 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_A6 = 1'b1;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_T1 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_B6 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_A1 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_A2 = CLBLM_R_X3Y6_SLICE_X2Y6_CQ;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_A3 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_A4 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_A5 = CLBLM_R_X3Y6_SLICE_X2Y6_C_XOR;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_A6 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_A1 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_AX = 1'b0;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_B1 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_B2 = CLBLM_R_X3Y6_SLICE_X2Y6_DQ;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_B3 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_B4 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_B5 = CLBLM_R_X3Y6_SLICE_X2Y6_D_XOR;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_B6 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_A3 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_A4 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_C6 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_BX = 1'b0;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_C1 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_C2 = CLBLM_R_X3Y6_SLICE_X2Y6_A_XOR;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_C3 = CLBLM_R_X3Y6_SLICE_X2Y6_AQ;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_C4 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_C5 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_C6 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_A5 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_A6 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_CIN = CLBLM_R_X3Y5_SLICE_X2Y5_COUT;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_CX = 1'b0;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_D1 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_D2 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_D3 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_D4 = CLBLM_R_X3Y6_SLICE_X2Y6_B_XOR;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_D5 = CLBLM_R_X3Y6_SLICE_X2Y6_BQ;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_D6 = 1'b1;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_DX = 1'b0;
  assign CLBLM_R_X3Y6_SLICE_X2Y6_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_B4 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_B5 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_B6 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_C5 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_C5 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_C6 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_A1 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_B1 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_A2 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_D1 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_A3 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_D2 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_D3 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_D1 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_D4 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_D2 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_D5 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_D6 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_A4 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_A5 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_A3 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_C6 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_A4 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_A5 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_A6 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_B1 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_A6 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_CX = 1'b0;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_A1 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_A2 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_A3 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_A4 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_A5 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_A6 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_A5 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_A6 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_B1 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_B2 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_B3 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_B4 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_B5 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_B6 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_B1 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_A1 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_B2 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_C1 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_C2 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_C3 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_C4 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_C5 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_C6 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_B3 = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_CE = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_B4 = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y8_CE = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_CE = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y11_CE = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_B5 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_D1 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_D2 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_D3 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_D4 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_D5 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X3Y7_D6 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_B6 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI15 = 1'b0;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_A1 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_A2 = CLBLL_L_X24Y46_SLICE_X36Y46_DQ;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_A3 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_A4 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_A5 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_A6 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_A4 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_A5 = CLBLM_R_X3Y7_SLICE_X2Y7_C_XOR;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_A6 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_A1 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_A2 = CLBLM_R_X3Y7_SLICE_X2Y7_CQ;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_AX = 1'b0;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_A3 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_B1 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_B2 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_B3 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_B4 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_B5 = CLBLM_R_X3Y7_SLICE_X2Y7_D_XOR;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_B1 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_B2 = CLBLM_R_X3Y7_SLICE_X2Y7_DQ;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_B3 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_B4 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_B5 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_B6 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_C1 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_C2 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_C4 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_C3 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_C4 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_C5 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_C6 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_CLK = RIOB33_X43Y25_IOB_X1Y26_I;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_C5 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_C6 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_CIN = CLBLM_R_X3Y6_SLICE_X2Y6_COUT;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_D1 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_D2 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_D3 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_D4 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_D5 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_D6 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_DX = CLBLL_L_X24Y46_SLICE_X36Y46_AO6;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_CX = 1'b0;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_D1 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_D2 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_D3 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_D4 = CLBLM_R_X3Y7_SLICE_X2Y7_B_XOR;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_D5 = CLBLM_R_X3Y7_SLICE_X2Y7_BQ;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_D6 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_DX = 1'b0;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_C6 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_C4 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_C5 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_A1 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_A2 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_A3 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_A4 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_A5 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_A6 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_B2 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_C6 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_B1 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_B2 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_B3 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_B4 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_B5 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_B6 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_D4 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_D5 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_D1 = LIOB33_X0Y5_IOB_X0Y6_I;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_C1 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_C2 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_C3 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_C4 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_C5 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_C6 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_D6 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y11_O;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_B1 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_D1 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_D1 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_D2 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_D3 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_D4 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_D5 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X37Y46_D6 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_D2 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_D3 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_D4 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_B2 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_D5 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_D1 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_A4 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_D6 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_D2 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_A2 = CLBLM_R_X11Y29_SLICE_X14Y29_CQ;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_D3 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_D4 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_B3 = 1'b1;
  assign LIOB33_X0Y43_IOB_X0Y43_O = CLBLM_R_X27Y43_SLICE_X43Y43_CQ;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_B4 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_B5 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_C5 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_C6 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_A1 = CLBLM_R_X27Y43_SLICE_X43Y43_C_XOR;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_B6 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_A2 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_A3 = CLBLM_R_X27Y38_SLICE_X43Y38_DQ;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_A4 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_A5 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_A6 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_AX = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_CIN = CLBLM_R_X27Y15_SLICE_X43Y15_COUT;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_B1 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_B2 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_B3 = CLBLM_R_X27Y41_SLICE_X43Y41_A5Q;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_B4 = CLBLM_R_X27Y43_SLICE_X43Y43_D_XOR;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_B5 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_B6 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_BX = 1'b0;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_B6 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_C1 = CLBLM_R_X27Y42_SLICE_X43Y42_A5Q;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_C2 = CLBLM_R_X27Y38_SLICE_X43Y38_D_XOR;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_BX = 1'b0;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_C3 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_C4 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_C5 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_C6 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_CX = 1'b0;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_D1 = CLBLM_R_X27Y38_SLICE_X43Y38_AO6;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_D2 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_D3 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_D4 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_D5 = CLBLM_R_X27Y38_SLICE_X43Y38_CQ;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_D6 = 1'b1;
  assign LIOB33_X0Y27_IOB_X0Y28_O = LIOB33_X0Y25_IOB_X0Y26_I;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_DX = 1'b0;
  assign CLBLM_R_X27Y38_SLICE_X43Y38_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_A1 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_A2 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_A3 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_A4 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_C5 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_A5 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_A6 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_B3 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_C6 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_B1 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_A1 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_A2 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_A3 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_A4 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_A5 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_A6 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_D3 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_D4 = CLBLM_R_X27Y16_SLICE_X43Y16_B_XOR;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_B2 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_B1 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_B2 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_B3 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_B4 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_B5 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_B6 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_CIN = CLBLM_R_X11Y28_SLICE_X14Y28_COUT;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_D5 = CLBLM_R_X27Y16_SLICE_X43Y16_BQ;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_C1 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_C2 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_C3 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_C4 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_C5 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_C6 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_D1 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_D2 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_D3 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_DX = 1'b0;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_D4 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_D5 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_D6 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_D1 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_D2 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_D3 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_D4 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_D5 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X3Y8_D6 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_A1 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_A2 = CLBLM_R_X3Y8_SLICE_X2Y8_AQ;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_A3 = CLBLM_R_X3Y9_SLICE_X2Y9_D_XOR;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_A4 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_A5 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_A6 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_A1 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_AX = 1'b0;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_B1 = CLBLM_R_X3Y8_SLICE_X2Y8_C_XOR;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_B2 = CLBLM_R_X3Y8_SLICE_X2Y8_DQ;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_B3 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_B4 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_B5 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_B6 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_A2 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_A3 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_A2 = CLBLM_R_X27Y42_SLICE_X43Y42_AQ;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_BX = 1'b0;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_D4 = CLBLM_R_X11Y29_SLICE_X14Y29_B_XOR;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_C1 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_C2 = CLBLM_R_X3Y8_SLICE_X2Y8_D_XOR;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_C3 = CLBLM_R_X3Y8_SLICE_X2Y8_BQ;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_C4 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_C5 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_C6 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_D5 = CLBLM_R_X11Y29_SLICE_X14Y29_BQ;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_A4 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_CIN = CLBLM_R_X3Y7_SLICE_X2Y7_COUT;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_A5 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_A6 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_A4 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_A5 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_CX = 1'b0;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_A6 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_D1 = CLBLM_R_X3Y8_SLICE_X2Y8_B_XOR;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_D2 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_D3 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_D4 = 1'b1;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_D5 = CLBLM_R_X3Y8_SLICE_X2Y8_CQ;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_D6 = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y11_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_O;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_DX = 1'b0;
  assign CLBLM_R_X3Y8_SLICE_X2Y8_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_AX = 1'b0;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_A6 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_B1 = CLBLM_R_X27Y42_SLICE_X43Y42_C_XOR;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_B1 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_T1 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_B2 = CLBLM_R_X27Y42_SLICE_X43Y42_DQ;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_B2 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_B3 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_B3 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_B4 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_B4 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_B5 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_B5 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_B6 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_C6 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_C1 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_C1 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_C2 = CLBLM_R_X27Y42_SLICE_X43Y42_D_XOR;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_CIN = CLBLM_R_X11Y5_SLICE_X15Y5_COUT;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_C2 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_C3 = CLBLM_R_X27Y42_SLICE_X43Y42_BQ;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O;
  assign LIOB33_X0Y17_IOB_X0Y18_O = CLBLM_R_X5Y20_SLICE_X7Y20_AQ;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_C3 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_C4 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DWE = 1'b0;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_C4 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_C5 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_C5 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_C6 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_C6 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_CIN = CLBLM_R_X27Y41_SLICE_X43Y41_COUT;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_D3 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_D4 = CLBLM_R_X11Y6_SLICE_X15Y6_B_XOR;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_CX = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSCLK = 1'b0;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_D5 = CLBLM_R_X11Y6_SLICE_X15Y6_BQ;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_D6 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_D1 = CLBLM_R_X27Y42_SLICE_X43Y42_B_XOR;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_D2 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_D3 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_D1 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_DX = 1'b0;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_D4 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_D2 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_A1 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_A2 = CLBLM_R_X27Y39_SLICE_X43Y39_CQ;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_D3 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_A3 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_A4 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_A5 = CLBLM_R_X27Y39_SLICE_X43Y39_C_XOR;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_A6 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_D4 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_AX = 1'b0;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_D5 = CLBLM_R_X27Y42_SLICE_X43Y42_CQ;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_B1 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_B2 = CLBLM_R_X27Y39_SLICE_X43Y39_DQ;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_B4 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_D5 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_B3 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_B4 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_B5 = CLBLM_R_X27Y39_SLICE_X43Y39_D_XOR;
  assign CLBLM_R_X27Y16_SLICE_X42Y16_D6 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_B6 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_BX = 1'b0;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_C1 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_C2 = CLBLM_R_X27Y39_SLICE_X43Y39_A_XOR;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_C3 = CLBLM_R_X27Y39_SLICE_X43Y39_AQ;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_C4 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_C5 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_C6 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_DX = 1'b0;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_CIN = CLBLM_R_X27Y38_SLICE_X43Y38_COUT;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSEN = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_CX = 1'b0;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_D1 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_D2 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_B5 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_A4 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_D3 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_D4 = CLBLM_R_X27Y39_SLICE_X43Y39_B_XOR;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_D5 = CLBLM_R_X27Y39_SLICE_X43Y39_BQ;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_D6 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_A6 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_A5 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_DX = 1'b0;
  assign CLBLM_R_X27Y39_SLICE_X43Y39_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_A1 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_A2 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_A3 = CLBLM_R_X5Y15_SLICE_X7Y15_DQ;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_A4 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_A5 = CLBLM_R_X5Y15_SLICE_X7Y15_C_XOR;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_A6 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_A6 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_A1 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_AX = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_A2 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_B1 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_B2 = CLBLM_R_X5Y15_SLICE_X7Y15_CQ;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_A1 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_B4 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_B5 = CLBLM_R_X5Y15_SLICE_X7Y15_D_XOR;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_B6 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_A2 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_A3 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_A4 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_A5 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_A6 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_BX = 1'b0;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_C4 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_C1 = CLBLM_R_X5Y15_SLICE_X7Y15_AQ;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_B1 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_B2 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_C5 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_C6 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_B3 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_B4 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_B5 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_B6 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_C1 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_C2 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_C3 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_C4 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_C5 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_C6 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_CX = 1'b0;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_D1 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_D2 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_D3 = CLBLM_R_X5Y15_SLICE_X7Y15_AO6;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_D4 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_D5 = CLBLM_R_X5Y15_SLICE_X7Y15_BQ;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_D6 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_DX = 1'b0;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_D1 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_D2 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_D3 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_D4 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_D5 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X3Y9_D6 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_A2 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_B1 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_B2 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_B3 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_A1 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_B4 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_B5 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_B6 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_A2 = CLBLM_R_X3Y9_SLICE_X2Y9_BQ;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_A3 = CLBLM_R_X3Y10_SLICE_X2Y10_D_XOR;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_A4 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_A5 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_C4 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_C5 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_C6 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_AX = 1'b0;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_B1 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_B2 = CLBLM_R_X3Y9_SLICE_X2Y9_DQ;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_B3 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_B4 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_B5 = CLBLM_R_X3Y9_SLICE_X2Y9_A_XOR;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_B6 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_BX = 1'b0;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_C1 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_C2 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_C3 = CLBLM_R_X3Y9_SLICE_X2Y9_CQ;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_C4 = CLBLM_R_X3Y10_SLICE_X2Y10_C_XOR;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_C5 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_D2 = 1'b1;
  assign CLBLL_L_X24Y46_SLICE_X36Y46_B6 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_D5 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_C6 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_D1 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_D6 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_CIN = CLBLM_R_X3Y8_SLICE_X2Y8_COUT;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_CX = 1'b0;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_D1 = CLBLM_R_X3Y9_SLICE_X2Y9_B_XOR;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_D2 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_D3 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_D4 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_D5 = CLBLM_R_X3Y8_SLICE_X2Y8_A5Q;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_D6 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_C4 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_C5 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_DX = 1'b0;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_C6 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_B3 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_C1 = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_CE = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_BX = CLBLL_L_X26Y9_SLICE_X40Y9_DQ;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_C2 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_C3 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_C3 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_C4 = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_CE = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_C5 = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_CE = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_C6 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_B4 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_C4 = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_CE = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_C4 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_D1 = 1'b1;
  assign LIOB33_X0Y19_IOB_X0Y19_O = CLBLM_R_X27Y19_SLICE_X43Y19_AQ;
  assign LIOB33_X0Y19_IOB_X0Y20_O = CLBLM_R_X11Y33_SLICE_X14Y33_AQ;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_D2 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_B5 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_D3 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_C5 = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_LOCKED;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_D4 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_C5 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_D5 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_D4 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_D6 = 1'b1;
  assign CLBLM_R_X3Y9_SLICE_X2Y9_A6 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_B6 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_C6 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_D1 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_D2 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_D3 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_D4 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_D5 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_BX = 1'b0;
  assign CLBLM_R_X27Y42_SLICE_X42Y42_D6 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_A1 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_A2 = CLBLM_R_X11Y32_SLICE_X14Y32_AQ;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_A3 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_A4 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_A5 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_CIN = CLBLM_R_X27Y18_SLICE_X43Y18_COUT;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_A6 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_AX = 1'b0;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_C1 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_A1 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_A1 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_A2 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_A3 = CLBLM_R_X27Y14_SLICE_X43Y14_DQ;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_B1 = CLBLM_R_X11Y32_SLICE_X14Y32_C_XOR;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_A4 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_A5 = CLBLM_R_X27Y14_SLICE_X43Y14_C_XOR;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_A6 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_A6 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_B2 = CLBLM_R_X11Y32_SLICE_X14Y32_DQ;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_AX = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_B1 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_B2 = CLBLM_R_X27Y14_SLICE_X43Y14_CQ;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_B3 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_B3 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_B4 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_B5 = CLBLM_R_X27Y14_SLICE_X43Y14_D_XOR;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_B6 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_C3 = CLBLM_R_X27Y19_SLICE_X43Y19_CQ;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_B4 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_C2 = CLBLM_R_X11Y32_SLICE_X14Y32_D_XOR;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_BX = 1'b0;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_C1 = CLBLM_R_X27Y14_SLICE_X43Y14_AQ;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_A1 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_A2 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_A3 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_A4 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_A5 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_A6 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_B5 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_B6 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_C3 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_B1 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_B2 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_B3 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_B4 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_B5 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_B6 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_CX = 1'b0;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_D1 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_D2 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_C1 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_C2 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_C3 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_C4 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_A1 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_A2 = CLBLM_R_X5Y16_SLICE_X7Y16_CQ;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_A3 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_A4 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_A5 = CLBLM_R_X5Y16_SLICE_X7Y16_C_XOR;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_A6 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_C5 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_C6 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_AX = 1'b0;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_B1 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_B2 = CLBLM_R_X5Y16_SLICE_X7Y16_DQ;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_A1 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_A2 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_B5 = CLBLM_R_X5Y16_SLICE_X7Y16_D_XOR;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_A3 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_B6 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_A4 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_A5 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_BX = 1'b0;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_C1 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_A6 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_C3 = CLBLM_R_X5Y16_SLICE_X7Y16_AQ;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_C2 = CLBLM_R_X5Y16_SLICE_X7Y16_A_XOR;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_A1 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_A2 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_A3 = CLBLM_R_X11Y28_SLICE_X14Y28_DQ;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_A4 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_A5 = CLBLM_R_X11Y28_SLICE_X14Y28_C_XOR;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_A6 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_C4 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_C5 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_C6 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_AX = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_CX = 1'b0;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_B1 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_B2 = CLBLM_R_X11Y28_SLICE_X14Y28_CQ;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_D1 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_D2 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_B3 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_D4 = CLBLM_R_X5Y16_SLICE_X7Y16_B_XOR;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_B4 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_B5 = CLBLM_R_X11Y28_SLICE_X14Y28_D_XOR;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_B6 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_BX = 1'b0;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_D5 = CLBLM_R_X5Y16_SLICE_X7Y16_BQ;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_C1 = CLBLM_R_X11Y28_SLICE_X14Y28_AQ;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_C2 = CLBLM_R_X11Y28_SLICE_X14Y28_B_XOR;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_C3 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_A2 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_C4 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_C5 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_C6 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X7Y16_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_D1 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_D2 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_D3 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_B1 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_B2 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_B3 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_CX = 1'b0;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_D1 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_D2 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_D3 = CLBLM_R_X11Y28_SLICE_X14Y28_AO6;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_D4 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_D5 = CLBLM_R_X11Y28_SLICE_X14Y28_BQ;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_D6 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_A1 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_C1 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_C2 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_DX = 1'b0;
  assign CLBLM_R_X11Y28_SLICE_X14Y28_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_AX = 1'b0;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_C3 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_C4 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_C5 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_C6 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_B1 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_B2 = CLBLM_R_X3Y10_SLICE_X2Y10_CQ;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_B3 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_B4 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_B5 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_B6 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_BX = 1'b0;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_C1 = CLBLM_R_X3Y10_SLICE_X2Y10_B_XOR;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_C2 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_C3 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_C4 = CLBLM_R_X3Y9_SLICE_X2Y9_C5Q;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_D3 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_D4 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_D5 = 1'b1;
  assign CLBLM_R_X5Y16_SLICE_X6Y16_D6 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_C6 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_CIN = CLBLM_R_X3Y9_SLICE_X2Y9_COUT;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_O;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_CX = 1'b0;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_D1 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_D2 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_D5 = CLBLM_R_X3Y9_SLICE_X2Y9_AQ;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_D6 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_D3 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_D4 = CLBLM_R_X3Y10_SLICE_X2Y10_A_XOR;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_DX = 1'b0;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_D3 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_D4 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_A3 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_A4 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_D5 = CLBLM_R_X11Y32_SLICE_X14Y32_CQ;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_D = LIOB33_X0Y11_IOB_X0Y12_I;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_A5 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_D6 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_A6 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_D1 = 1'b1;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_D = LIOB33_X0Y11_IOB_X0Y11_I;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_DX = 1'b0;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_CIN = CLBLM_R_X11Y31_SLICE_X14Y31_COUT;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_B1 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_D2 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_B2 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_B3 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_B4 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_B5 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_B6 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_D3 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_D4 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_DX = 1'b0;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_C1 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_C2 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_C3 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_C4 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_C5 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_C2 = CLBLM_R_X27Y14_SLICE_X43Y14_B_XOR;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_D5 = CLBLM_R_X27Y19_SLICE_X43Y19_DQ;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_C6 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_C4 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_C5 = 1'b1;
  assign LIOI3_X0Y27_OLOGIC_X0Y28_D1 = LIOB33_X0Y25_IOB_X0Y26_I;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_C6 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_C5 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_D6 = 1'b1;
  assign LIOI3_X0Y27_OLOGIC_X0Y28_T1 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_C3 = CLBLM_R_X11Y31_SLICE_X14Y31_BQ;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_A1 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_A2 = CLBLM_R_X27Y41_SLICE_X43Y41_AQ;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_A1 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_A2 = CLBLM_R_X27Y15_SLICE_X43Y15_CQ;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_A3 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_A4 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_A5 = CLBLM_R_X27Y15_SLICE_X43Y15_C_XOR;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_A6 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_A3 = CLBLM_R_X27Y38_SLICE_X43Y38_B_XOR;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_A4 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_AX = 1'b0;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_B1 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_B2 = CLBLM_R_X27Y15_SLICE_X43Y15_DQ;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_B3 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_B4 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_B5 = CLBLM_R_X27Y15_SLICE_X43Y15_D_XOR;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_B6 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_B1 = CLBLM_R_X27Y41_SLICE_X43Y41_C_XOR;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_B2 = CLBLM_R_X27Y41_SLICE_X43Y41_DQ;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_BX = 1'b0;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_D1 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_C1 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_C4 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_A1 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_A2 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_A3 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_A4 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_A5 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_A6 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_C2 = CLBLM_R_X27Y15_SLICE_X43Y15_A_XOR;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_CX = 1'b0;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_C3 = CLBLM_R_X27Y15_SLICE_X43Y15_AQ;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_B1 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_B2 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_B3 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_B4 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_B5 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_B6 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_CX = 1'b0;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_D1 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_D3 = CLBLM_R_X27Y14_SLICE_X43Y14_AO6;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_C1 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_C2 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_C3 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_C4 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_A1 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_A2 = CLBLM_R_X5Y17_SLICE_X7Y17_CQ;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_A3 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_A4 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_A5 = CLBLM_R_X5Y17_SLICE_X7Y17_C_XOR;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_A6 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_C5 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_C6 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_AX = 1'b0;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_B1 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_B2 = CLBLM_R_X5Y17_SLICE_X7Y17_DQ;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_B3 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_B4 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_B5 = CLBLM_R_X5Y17_SLICE_X7Y17_D_XOR;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_B6 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_D1 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_D2 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_BX = 1'b0;
  assign CLBLM_R_X11Y29_SLICE_X15Y29_D3 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_C1 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_C2 = CLBLM_R_X5Y17_SLICE_X7Y17_A_XOR;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_C3 = CLBLM_R_X5Y17_SLICE_X7Y17_AQ;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_C4 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_C5 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_C6 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_A3 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_CIN = CLBLM_R_X5Y16_SLICE_X7Y16_COUT;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_A4 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_A5 = CLBLM_R_X11Y29_SLICE_X14Y29_C_XOR;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_A6 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_A1 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_CX = 1'b0;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_AX = 1'b0;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_D1 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_D2 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_D3 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_D4 = CLBLM_R_X5Y17_SLICE_X7Y17_B_XOR;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_D5 = CLBLM_R_X5Y17_SLICE_X7Y17_BQ;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_D6 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_B1 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_B2 = CLBLM_R_X11Y29_SLICE_X14Y29_DQ;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_DX = 1'b0;
  assign CLBLM_R_X5Y17_SLICE_X7Y17_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_B3 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_B4 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_B5 = CLBLM_R_X11Y29_SLICE_X14Y29_D_XOR;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_A1 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_A2 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_A3 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_A4 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_A5 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_A6 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_C1 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_C2 = CLBLM_R_X11Y29_SLICE_X14Y29_A_XOR;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_C3 = CLBLM_R_X11Y29_SLICE_X14Y29_AQ;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_C4 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_B1 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_B2 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_B3 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_B4 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_B5 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_B6 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_CX = 1'b0;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_D1 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_D2 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_D3 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_C1 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_C2 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_C3 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_C4 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_C5 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_C6 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_D6 = 1'b1;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_DX = 1'b0;
  assign CLBLM_R_X11Y29_SLICE_X14Y29_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_A6 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_CX = 1'b0;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_D1 = CLBLM_R_X27Y18_SLICE_X43Y18_B_XOR;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_A5 = CLBLM_R_X27Y40_SLICE_X43Y40_C_XOR;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_D1 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_D2 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_D3 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_D4 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_D5 = 1'b1;
  assign CLBLM_R_X5Y17_SLICE_X6Y17_D6 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_AX = 1'b0;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_CIN = CLBLM_R_X11Y30_SLICE_X14Y30_COUT;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_D1 = CLBLM_R_X11Y32_SLICE_X14Y32_B_XOR;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_D2 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_B1 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_B1 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_B2 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_B2 = CLBLM_R_X27Y40_SLICE_X43Y40_DQ;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_B3 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_B3 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_B4 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_B4 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_B5 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_B5 = CLBLM_R_X27Y40_SLICE_X43Y40_D_XOR;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_D3 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_B6 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_B6 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_A1 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_BX = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR0 = 1'b0;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_D = LIOB33_X0Y9_IOB_X0Y10_I;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR1 = 1'b0;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_D4 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_C1 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR2 = 1'b0;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_C2 = CLBLM_R_X27Y40_SLICE_X43Y40_A_XOR;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_C1 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR3 = 1'b0;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_A2 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_C3 = CLBLM_R_X27Y40_SLICE_X43Y40_AQ;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_C2 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR4 = 1'b0;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_C4 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_C3 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR5 = 1'b0;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_C5 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_C4 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR6 = 1'b0;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_D5 = CLBLM_R_X27Y18_SLICE_X43Y18_CQ;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_C6 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_C5 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DCLK = 1'b0;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_C6 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DEN = 1'b0;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_CIN = CLBLM_R_X27Y39_SLICE_X43Y39_COUT;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI0 = 1'b0;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI1 = 1'b0;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_C6 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI2 = 1'b0;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_D6 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI3 = 1'b0;
  assign LIOB33_SING_X0Y0_IOB_X0Y0_O = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_LOCKED;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI4 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI5 = 1'b0;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_CX = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI6 = 1'b0;
  assign CLBLM_R_X11Y32_SLICE_X14Y32_D2 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI7 = 1'b0;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_D1 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI8 = 1'b0;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_D2 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI9 = 1'b0;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_D1 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_D3 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI10 = 1'b0;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_D2 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_D4 = CLBLM_R_X27Y40_SLICE_X43Y40_B_XOR;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI11 = 1'b0;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_D3 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_D5 = CLBLM_R_X27Y40_SLICE_X43Y40_BQ;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI12 = 1'b0;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_D4 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_D6 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI13 = 1'b0;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_D5 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI14 = 1'b0;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_D6 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_C5 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_A1 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_A1 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_A2 = CLBLM_R_X27Y16_SLICE_X43Y16_CQ;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_A3 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_A4 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_A5 = CLBLM_R_X27Y16_SLICE_X43Y16_C_XOR;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_A6 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_DX = 1'b0;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_AX = 1'b0;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_DX = 1'b0;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_B1 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_B2 = CLBLM_R_X27Y16_SLICE_X43Y16_DQ;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_B3 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_B4 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_B5 = CLBLM_R_X27Y16_SLICE_X43Y16_D_XOR;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_B6 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_B6 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_BX = 1'b0;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_BX = 1'b0;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_C1 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_C2 = CLBLM_R_X27Y16_SLICE_X43Y16_A_XOR;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_A1 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_C6 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_A2 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_A3 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_A4 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_A5 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_A6 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_C3 = CLBLM_R_X27Y16_SLICE_X43Y16_AQ;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_C4 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_B1 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_B2 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_B3 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_B4 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_B5 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_B6 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_CX = 1'b0;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_D1 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_D2 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_C1 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_C2 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_C3 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_C4 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_A1 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_A2 = CLBLM_R_X5Y18_SLICE_X7Y18_AQ;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_A3 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_A4 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_A5 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_A6 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_C5 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_C6 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_AX = 1'b0;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_B1 = CLBLM_R_X5Y18_SLICE_X7Y18_C_XOR;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_B2 = CLBLM_R_X5Y18_SLICE_X7Y18_DQ;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_B3 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_B4 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_B5 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_B6 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_D1 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_D2 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_BX = 1'b0;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_D3 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_C1 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_C2 = CLBLM_R_X5Y18_SLICE_X7Y18_D_XOR;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_C3 = CLBLM_R_X5Y18_SLICE_X7Y18_BQ;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_C4 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_C5 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_C6 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_A1 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_CIN = CLBLM_R_X5Y17_SLICE_X7Y17_COUT;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_A2 = CLBLM_R_X11Y30_SLICE_X14Y30_CQ;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_A3 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_A4 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_A5 = CLBLM_R_X11Y30_SLICE_X14Y30_C_XOR;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_CX = 1'b0;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_A6 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_D1 = CLBLM_R_X5Y18_SLICE_X7Y18_B_XOR;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_D2 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_D3 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_D4 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_D5 = CLBLM_R_X5Y18_SLICE_X7Y18_CQ;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_D6 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_AX = 1'b0;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_B1 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_DX = 1'b0;
  assign CLBLM_R_X5Y18_SLICE_X7Y18_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_B2 = CLBLM_R_X11Y30_SLICE_X14Y30_DQ;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_B3 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_B4 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_A1 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_A2 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_A3 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_A4 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_A5 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_A6 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_C1 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_C2 = CLBLM_R_X11Y30_SLICE_X14Y30_A_XOR;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_C3 = CLBLM_R_X11Y30_SLICE_X14Y30_AQ;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_C4 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_B1 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_B2 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_B3 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_B4 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_B5 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_B6 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_CX = 1'b0;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_D1 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_D2 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_D3 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_C1 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_C2 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_C3 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_C4 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_C5 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_C6 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_D6 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_DX = 1'b0;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_D3 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_RST = CLBLM_R_X27Y8_SLICE_X42Y8_DQ;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_D1 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_D2 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_D3 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_D4 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_D5 = 1'b1;
  assign CLBLM_R_X5Y18_SLICE_X6Y18_D6 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_C1 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_C2 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_C3 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_D4 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_C4 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_C5 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_C6 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_D5 = CLBLM_R_X27Y17_SLICE_X43Y17_CQ;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_D4 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_D5 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_D6 = 1'b1;
  assign RIOI3_X43Y25_ILOGIC_X1Y26_D = RIOB33_X43Y25_IOB_X1Y26_I;
  assign CLBLM_R_X11Y30_SLICE_X15Y30_D6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_T1 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_D1 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_D2 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_D3 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_D4 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_D5 = 1'b1;
  assign CLBLM_R_X27Y40_SLICE_X42Y40_D6 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_DX = 1'b0;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_BX = 1'b0;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_C1 = 1'b1;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_C2 = CLBLM_R_X3Y7_SLICE_X2Y7_A_XOR;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X3Y7_SLICE_X2Y7_C3 = CLBLM_R_X3Y7_SLICE_X2Y7_AQ;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_B6 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_C3 = CLBLM_R_X27Y17_SLICE_X43Y17_BQ;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_C4 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_A1 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_A1 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_A2 = CLBLM_R_X27Y17_SLICE_X43Y17_AQ;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_A3 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_A4 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_A5 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_B5 = CLBLM_R_X11Y30_SLICE_X14Y30_D_XOR;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_A6 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_C5 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_AX = 1'b0;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_C6 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_B6 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_B1 = CLBLM_R_X27Y17_SLICE_X43Y17_C_XOR;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_B2 = CLBLM_R_X27Y17_SLICE_X43Y17_DQ;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_B3 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_B4 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_B5 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_B6 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_B1 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_BX = 1'b0;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_CIN = CLBLM_R_X27Y16_SLICE_X43Y16_COUT;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_C1 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_C2 = CLBLM_R_X27Y17_SLICE_X43Y17_D_XOR;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_A1 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_A2 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_A1 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_A2 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_A3 = CLBLM_R_X11Y5_SLICE_X15Y5_DQ;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_A4 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_A5 = CLBLM_R_X11Y5_SLICE_X15Y5_C_XOR;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_A6 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_BX = 1'b0;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_A3 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_AX = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_A4 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_B1 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_B2 = CLBLM_R_X11Y5_SLICE_X15Y5_CQ;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_B3 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_B4 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_B5 = CLBLM_R_X11Y5_SLICE_X15Y5_D_XOR;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_B6 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_B1 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_B2 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_BX = 1'b0;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_B3 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_C1 = CLBLM_R_X11Y5_SLICE_X15Y5_AQ;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_C2 = CLBLM_R_X11Y5_SLICE_X15Y5_B_XOR;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_A1 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_A2 = CLBLM_R_X5Y19_SLICE_X7Y19_AQ;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_A3 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_A4 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_A5 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_A6 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_C3 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_C4 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_AX = 1'b0;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_C5 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_B1 = CLBLM_R_X5Y19_SLICE_X7Y19_C_XOR;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_B2 = CLBLM_R_X5Y19_SLICE_X7Y19_DQ;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_B3 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_B4 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_B5 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_B6 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_CX = 1'b0;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_D1 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_BX = 1'b0;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_D2 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_C1 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_DX = 1'b0;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_C2 = CLBLM_R_X5Y19_SLICE_X7Y19_D_XOR;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_C3 = CLBLM_R_X5Y19_SLICE_X7Y19_BQ;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_C4 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_C5 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_C6 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_CIN = CLBLM_R_X5Y18_SLICE_X7Y18_COUT;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_A1 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_A2 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_A3 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_A4 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_CX = 1'b0;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_A5 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_D1 = CLBLM_R_X5Y19_SLICE_X7Y19_B_XOR;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_D2 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_D3 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_D4 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_D5 = CLBLM_R_X5Y19_SLICE_X7Y19_CQ;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_D6 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_B1 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_B2 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_DX = 1'b0;
  assign CLBLM_R_X5Y19_SLICE_X7Y19_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_B3 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_B4 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_B5 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_A1 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_A2 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_A3 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_A4 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_A5 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_A6 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_C1 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_C2 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_C3 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_B1 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_B2 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_B3 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_B4 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_B5 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_B6 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_D1 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_D2 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_D3 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_C1 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_C2 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_C3 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_C4 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_C5 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_C6 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_D4 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_D5 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_D6 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_DX = 1'b0;
  assign CLBLM_R_X11Y31_SLICE_X14Y31_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_A1 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_A2 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_D1 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_D2 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_D3 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_D4 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_D5 = 1'b1;
  assign CLBLM_R_X5Y19_SLICE_X6Y19_D6 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_D4 = CLBLM_R_X11Y30_SLICE_X14Y30_B_XOR;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_A3 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_A4 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_D5 = CLBLM_R_X11Y30_SLICE_X14Y30_BQ;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_A3 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_A5 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_A2 = CLBLM_R_X27Y43_SLICE_X43Y43_DQ;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_A4 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_A5 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_A6 = 1'b1;
  assign CLBLM_R_X27Y16_SLICE_X43Y16_D6 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_A6 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_AX = 1'b0;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_B1 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_B2 = CLBLM_R_X27Y43_SLICE_X43Y43_CQ;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_B2 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_B3 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_B3 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_B4 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_B4 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_B5 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_B5 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_B6 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_B6 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_BX = 1'b0;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_C1 = CLBLM_R_X27Y43_SLICE_X43Y43_B_XOR;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_B3 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_C1 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_C2 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_C2 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_C3 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_C3 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_C4 = CLBLM_R_X27Y38_SLICE_X43Y38_AQ;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_C4 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_C5 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_C5 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_C6 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_C6 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_CIN = CLBLM_R_X27Y42_SLICE_X43Y42_COUT;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_C2 = CLBLM_R_X5Y15_SLICE_X7Y15_B_XOR;
  assign CLBLM_R_X5Y15_SLICE_X7Y15_C3 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PWRDWN = LIOB33_X0Y11_IOB_X0Y12_I;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_CX = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBIN = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBOUT;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKIN1 = CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y8_O;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_D1 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSINCDEC = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKIN2 = RIOB33_X43Y25_IOB_X1Y26_I;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKINSEL = LIOB33_X0Y9_IOB_X0Y10_I;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_D2 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_D3 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_D1 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_A1 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_A2 = CLBLM_R_X27Y18_SLICE_X43Y18_AQ;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_A3 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_A4 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_D2 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_A5 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_A6 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_AX = 1'b0;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_D3 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_B1 = CLBLM_R_X27Y18_SLICE_X43Y18_C_XOR;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_B2 = CLBLM_R_X27Y18_SLICE_X43Y18_DQ;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_B3 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_B4 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_D4 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_B5 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_B6 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_BX = 1'b0;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_B1 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_D5 = 1'b1;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_C1 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_A1 = 1'b1;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_A2 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_A1 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_A2 = CLBLM_R_X11Y6_SLICE_X15Y6_CQ;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_A3 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_A4 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_A5 = CLBLM_R_X11Y6_SLICE_X15Y6_C_XOR;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_A6 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_B2 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_B3 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_AX = 1'b0;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_A3 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_B1 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_B2 = CLBLM_R_X11Y6_SLICE_X15Y6_DQ;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_B3 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_B4 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_B5 = CLBLM_R_X11Y6_SLICE_X15Y6_D_XOR;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_B6 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_B4 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_B5 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_BX = 1'b0;
  assign CLBLM_R_X11Y32_SLICE_X15Y32_B3 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_C1 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_C2 = CLBLM_R_X11Y6_SLICE_X15Y6_A_XOR;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_A1 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_A2 = CLBLM_R_X5Y20_SLICE_X7Y20_BQ;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_A3 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_A4 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_A5 = CLBLM_R_X5Y20_SLICE_X7Y20_B_XOR;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_A6 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_C3 = CLBLM_R_X11Y6_SLICE_X15Y6_AQ;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_C4 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_AX = 1'b0;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_C5 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_B1 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_B2 = CLBLM_R_X5Y20_SLICE_X7Y20_AQ;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_B3 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_B4 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_B5 = CLBLM_R_X5Y20_SLICE_X7Y20_A_XOR;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_B6 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_CX = 1'b0;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_D1 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_BX = 1'b0;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_D2 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_C1 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_C2 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_C3 = CLBLM_R_X5Y20_SLICE_X7Y20_CQ;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_C4 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_C5 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_C6 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_A1 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_CIN = CLBLM_R_X5Y19_SLICE_X7Y19_COUT;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_O;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_A2 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_A3 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X15Y6_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_A4 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_CX = 1'b0;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_A5 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_D1 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_D2 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_D3 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_D4 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_D5 = CLBLM_R_X5Y20_SLICE_X7Y20_DQ;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_D6 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_B5 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_B6 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_B1 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_DX = 1'b0;
  assign CLBLM_R_X5Y20_SLICE_X7Y20_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_B2 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_B3 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_B4 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_A1 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_A2 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_A3 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_A4 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_A5 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_A6 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_C1 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_C2 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_C3 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_B1 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_B2 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_B3 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_B4 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_B5 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_B6 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_D1 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_D2 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_D3 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_C1 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_C2 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_C3 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_C4 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_C5 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_C6 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_D5 = 1'b1;
  assign CLBLM_R_X11Y6_SLICE_X14Y6_D6 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_A5 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_A6 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_A3 = CLBLM_R_X27Y38_SLICE_X43Y38_C_XOR;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_B4 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_D1 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_D2 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_D3 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_D4 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_D5 = 1'b1;
  assign CLBLM_R_X5Y20_SLICE_X6Y20_D6 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_C2 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_B5 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_B6 = 1'b1;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_D1 = CLBLM_R_X5Y20_SLICE_X7Y20_AQ;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_D4 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_A1 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_A2 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_A3 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_A4 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_A5 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_A6 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_D5 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_C1 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_D6 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_B1 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_B2 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_B3 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_B4 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_B5 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_B6 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_C2 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_C3 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_C1 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_C2 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_C3 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_C4 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_C5 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_C6 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_C4 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y11_O;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_C5 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_C6 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_D1 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_D2 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_D3 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_D4 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_D5 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_D6 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X40Y9_DX = LIOB33_X0Y11_IOB_X0Y11_I;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_C1 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_A2 = CLBLM_R_X3Y10_SLICE_X2Y10_DQ;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_C2 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_D3 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_D2 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_A3 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_C3 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_A4 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_D5 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_A1 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_A2 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_A3 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_A4 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_A5 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_A6 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_A5 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_A6 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_D6 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_B1 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_B2 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_B3 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_B4 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_B5 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_B6 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_D3 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_D1 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_C1 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_C2 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_C3 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_C4 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_C5 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_C6 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_D2 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_D3 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_D4 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_D1 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_D2 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_D3 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_D4 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_D5 = 1'b1;
  assign CLBLL_L_X26Y9_SLICE_X41Y9_D6 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_D4 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_D5 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_D6 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_D5 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_D3 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_D4 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_A1 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_A2 = CLBLM_R_X27Y19_SLICE_X43Y19_BQ;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_A3 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_AX = 1'b0;
  assign CLBLM_R_X27Y19_SLICE_X42Y19_D6 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_A4 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_A5 = CLBLM_R_X27Y19_SLICE_X43Y19_B_XOR;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_A6 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_AX = 1'b0;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_B1 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_D4 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_B2 = CLBLM_R_X27Y19_SLICE_X43Y19_AQ;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_B3 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_B4 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_B5 = CLBLM_R_X27Y19_SLICE_X43Y19_A_XOR;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_B6 = 1'b1;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_C1 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_BX = 1'b0;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_C1 = 1'b1;
  assign CLBLM_R_X27Y19_SLICE_X43Y19_C2 = CLBLM_R_X27Y8_SLICE_X42Y8_DQ;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_A1 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_A2 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_A1 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_A2 = CLBLM_R_X11Y7_SLICE_X15Y7_CQ;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_A3 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_A4 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_A5 = CLBLM_R_X11Y7_SLICE_X15Y7_C_XOR;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_A6 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X2Y10_C5 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_B4 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_AX = 1'b0;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_B5 = CLBLM_R_X11Y33_SLICE_X14Y33_A_XOR;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_B1 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_B2 = CLBLM_R_X11Y7_SLICE_X15Y7_DQ;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_B3 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_B4 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_B5 = CLBLM_R_X11Y7_SLICE_X15Y7_D_XOR;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_B6 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_B6 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_B1 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_BX = 1'b0;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_B3 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_C1 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_C2 = CLBLM_R_X11Y7_SLICE_X15Y7_A_XOR;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_C3 = CLBLM_R_X11Y7_SLICE_X15Y7_AQ;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_C4 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_C5 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_C6 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_C1 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_CIN = CLBLM_R_X11Y6_SLICE_X15Y6_COUT;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_C3 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_C4 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_C5 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_C6 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_CX = 1'b0;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_BX = 1'b0;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_D1 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_D2 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_D3 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_D4 = CLBLM_R_X11Y7_SLICE_X15Y7_B_XOR;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_D5 = CLBLM_R_X11Y7_SLICE_X15Y7_BQ;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_D6 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_D1 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_D2 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_DX = 1'b0;
  assign CLBLM_R_X11Y7_SLICE_X15Y7_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_D4 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_A1 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_A2 = CLBLM_R_X11Y33_SLICE_X14Y33_BQ;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_A1 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_A2 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_A3 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_A4 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_A5 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_A6 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_A3 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_A4 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_A5 = CLBLM_R_X11Y33_SLICE_X14Y33_B_XOR;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_A6 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_B1 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_B2 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_B3 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_B4 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_B5 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_B6 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_B1 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_B2 = CLBLM_R_X11Y33_SLICE_X14Y33_AQ;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_B3 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_C1 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_C1 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_C2 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_C3 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_C4 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_C5 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_C6 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_C2 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_C3 = CLBLM_R_X11Y33_SLICE_X14Y33_CQ;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_C4 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_C5 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_C6 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_CIN = CLBLM_R_X11Y32_SLICE_X14Y32_COUT;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_O;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_CX = 1'b0;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_D1 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_D1 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_D2 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_D3 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_D4 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_D5 = 1'b1;
  assign CLBLM_R_X11Y7_SLICE_X14Y7_D6 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_D2 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_D3 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_D4 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_D5 = CLBLM_R_X11Y33_SLICE_X14Y33_DQ;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_D6 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_DX = 1'b0;
  assign CLBLM_R_X11Y33_SLICE_X14Y33_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_C1 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_C2 = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y0_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_O;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_C3 = 1'b1;
  assign LIOB33_X0Y3_IOB_X0Y4_O = CLBLM_R_X11Y10_SLICE_X15Y10_AQ;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_C4 = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y3_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_O;
  assign LIOB33_X0Y3_IOB_X0Y3_O = CLBLM_R_X3Y10_SLICE_X2Y10_CQ;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_DX = 1'b0;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_C5 = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_O;
  assign CLBLM_R_X27Y39_SLICE_X42Y39_C2 = 1'b1;
  assign CLBLM_R_X27Y38_SLICE_X42Y38_C6 = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y6_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_D1 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X43Y14_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_D2 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_D3 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_D4 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_D5 = 1'b1;
  assign CLBLM_R_X11Y28_SLICE_X15Y28_D6 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_A2 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_CX = 1'b0;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_D1 = CLBLM_R_X11Y10_SLICE_X15Y10_AQ;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_O;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y8_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_O;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_T1 = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_D1 = CLBLM_R_X3Y10_SLICE_X2Y10_CQ;
  assign CLBLM_R_X27Y18_SLICE_X43Y18_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_T1 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_A1 = 1'b1;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_T1 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_A2 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_C4 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_C5 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_C6 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_A3 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_CIN = CLBLM_R_X27Y14_SLICE_X43Y14_COUT;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_A2 = CLBLM_R_X27Y40_SLICE_X43Y40_CQ;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y7_O;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_D4 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_D5 = CLBLM_R_X11Y10_SLICE_X15Y10_DQ;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_D6 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_A4 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_A1 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_A2 = CLBLM_R_X11Y8_SLICE_X15Y8_AQ;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_A3 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_A4 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_A5 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_A6 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_DX = 1'b0;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_A3 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_AX = 1'b0;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_B1 = CLBLM_R_X11Y8_SLICE_X15Y8_C_XOR;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_B2 = CLBLM_R_X11Y8_SLICE_X15Y8_DQ;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_B3 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_B4 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_B5 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_B6 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X15Y10_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_BX = 1'b0;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_C1 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_C2 = CLBLM_R_X11Y8_SLICE_X15Y8_D_XOR;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_C3 = CLBLM_R_X11Y8_SLICE_X15Y8_BQ;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_C4 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_C5 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_C6 = 1'b1;
  assign CLBLM_R_X27Y14_SLICE_X42Y14_A5 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_CIN = CLBLM_R_X11Y7_SLICE_X15Y7_COUT;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_D2 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_D3 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_D4 = CLBLM_R_X27Y15_SLICE_X43Y15_B_XOR;
  assign CLBLM_R_X27Y40_SLICE_X43Y40_A4 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_CX = 1'b0;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_D1 = CLBLM_R_X11Y8_SLICE_X15Y8_B_XOR;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_D2 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_D3 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_D4 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_D5 = CLBLM_R_X11Y8_SLICE_X15Y8_CQ;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_D6 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_D5 = CLBLM_R_X27Y15_SLICE_X43Y15_BQ;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_D6 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_DX = 1'b0;
  assign CLBLM_R_X11Y8_SLICE_X15Y8_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_A4 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_A1 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_A2 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_A3 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_A4 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_A5 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_A6 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_DX = 1'b0;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_B1 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_B2 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_B3 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_B4 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_B5 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_B6 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_B6 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X43Y15_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_C1 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_C2 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_C3 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_C4 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_C5 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_C6 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_A1 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_D1 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_D2 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_D3 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_D4 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_D5 = 1'b1;
  assign CLBLM_R_X11Y8_SLICE_X14Y8_D6 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_A2 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_A3 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_A4 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_A5 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_A5 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_A6 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_D4 = CLBLM_R_X27Y43_SLICE_X43Y43_A_XOR;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_D1 = CLBLM_R_X27Y17_SLICE_X43Y17_B_XOR;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_A6 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_B6 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_AX = 1'b0;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_D5 = CLBLM_R_X27Y38_SLICE_X43Y38_BQ;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_B1 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_B2 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_B3 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_B3 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_B4 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_B4 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_D6 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_B5 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_B5 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_B6 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_B6 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_C6 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_BX = 1'b0;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_C6 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_C1 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_C1 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_C1 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_C2 = CLBLM_R_X27Y41_SLICE_X43Y41_D_XOR;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_A3 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_C2 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_C3 = CLBLM_R_X27Y41_SLICE_X43Y41_BQ;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_C4 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_C3 = 1'b1;
  assign CLBLM_R_X27Y17_SLICE_X42Y17_D6 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_C5 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_C4 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_C6 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_C5 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_C2 = 1'b1;
  assign CLBLM_R_X11Y30_SLICE_X14Y30_CIN = CLBLM_R_X11Y29_SLICE_X14Y29_COUT;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_C6 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_A4 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_CIN = CLBLM_R_X27Y40_SLICE_X43Y40_COUT;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X1Y10_O;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_DX = 1'b0;
  assign CLBLM_R_X27Y17_SLICE_X43Y17_D2 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_D4 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_C3 = 1'b1;
  assign CLBLM_R_X11Y10_SLICE_X14Y10_D5 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_D3 = CLBLM_R_X11Y5_SLICE_X15Y5_AO6;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_A5 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_D4 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_CX = 1'b0;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_D5 = CLBLM_R_X11Y5_SLICE_X15Y5_BQ;
  assign CLBLM_R_X27Y43_SLICE_X43Y43_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_D6 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_D1 = CLBLM_R_X27Y41_SLICE_X43Y41_B_XOR;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_C4 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_D2 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_A6 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_D3 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_D1 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_D4 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_D2 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X15Y5_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1 = CLBLM_R_X27Y43_SLICE_X43Y43_CQ;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_D5 = CLBLM_R_X27Y41_SLICE_X43Y41_CQ;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_D3 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_D6 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_D4 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_C5 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_A1 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_A2 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_A3 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_A4 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_A5 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_A6 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_D5 = 1'b1;
  assign CLBLM_R_X27Y15_SLICE_X42Y15_D6 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_B1 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_B2 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_B3 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_B4 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_B5 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_B6 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_DX = 1'b0;
  assign CLBLM_R_X27Y41_SLICE_X43Y41_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_C1 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_C2 = 1'b1;
  assign CLBLM_R_X3Y10_SLICE_X3Y10_C6 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_A1 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_A2 = CLBLM_R_X11Y9_SLICE_X15Y9_AQ;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_A3 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_A4 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_A5 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_A6 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_C3 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X43Y8_C4 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_AX = 1'b0;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_A6 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_B1 = CLBLM_R_X11Y9_SLICE_X15Y9_C_XOR;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_B2 = CLBLM_R_X11Y9_SLICE_X15Y9_DQ;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_B3 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_B4 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_B5 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_B6 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_A5 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_A6 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_BX = 1'b0;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_C1 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_C2 = CLBLM_R_X11Y9_SLICE_X15Y9_D_XOR;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_C3 = CLBLM_R_X11Y9_SLICE_X15Y9_BQ;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_C4 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_C5 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_C6 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_A1 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_CIN = CLBLM_R_X11Y8_SLICE_X15Y8_COUT;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y4_O;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_A2 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_A3 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_CX = 1'b0;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_A4 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_D1 = CLBLM_R_X11Y9_SLICE_X15Y9_B_XOR;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_D2 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_D3 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_D4 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_D5 = CLBLM_R_X11Y9_SLICE_X15Y9_CQ;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_D6 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_DX = 1'b0;
  assign CLBLM_R_X11Y9_SLICE_X15Y9_SR = CLBLM_R_X27Y19_SLICE_X43Y19_CO5;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_B1 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_B2 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_B3 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_A1 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_A2 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_A3 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_A4 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_A5 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_A6 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_B4 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_C1 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_C2 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_C3 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_B1 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_B2 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_B3 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_B4 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_B5 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_B6 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_B6 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_B5 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_B6 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_CX = CLBLM_R_X27Y8_SLICE_X42Y8_BQ;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_C1 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_C2 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_C3 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_C4 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_C5 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_C6 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_D5 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_D6 = 1'b1;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_DX = CLBLM_R_X27Y8_SLICE_X42Y8_CQ;
  assign CLBLM_R_X27Y8_SLICE_X42Y8_SR = LIOB33_X0Y11_IOB_X0Y11_I;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_B2 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_A1 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_B3 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_B4 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_D1 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_D2 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_D3 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_D4 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_D5 = 1'b1;
  assign CLBLM_R_X11Y9_SLICE_X14Y9_D6 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_C1 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_B5 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_C2 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_B6 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_A3 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_C3 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_C4 = 1'b1;
  assign CLBLM_R_X27Y42_SLICE_X43Y42_D6 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_C5 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_C4 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_B2 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_C6 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_C5 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_A4 = 1'b1;
  assign CLBLM_R_X11Y5_SLICE_X14Y5_C6 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_C1 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_C2 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0 = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT0;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_A3 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_C3 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I0 = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I1 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_C4 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_C5 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_A5 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_C6 = 1'b1;
  assign CLBLM_R_X5Y15_SLICE_X6Y15_A4 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_B4 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_I0 = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT2;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_I1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_I0 = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT3;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_I1 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_D1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_I0 = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT4;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y12_I1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_I0 = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT5;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_D2 = 1'b1;
  assign CLBLM_R_X27Y43_SLICE_X42Y43_A6 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y13_I1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_I0 = RIOB33_X43Y25_IOB_X1Y26_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y14_I1 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_D3 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_I0 = RIOB33_X43Y25_IOB_X1Y26_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y15_I1 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_D4 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_D5 = 1'b1;
  assign CLBLM_R_X11Y33_SLICE_X15Y33_B5 = 1'b1;
  assign CLBLM_R_X11Y31_SLICE_X15Y31_D6 = 1'b1;
  assign CLBLM_R_X27Y41_SLICE_X42Y41_D1 = 1'b1;
endmodule
