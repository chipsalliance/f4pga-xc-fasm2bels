module top(
  input clk,
  input jc1,
  input jc3,
  input [7:0] sw,
  output jc2,
  output jc4,
  output [7:0] led
  );
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_A;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_A1;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_A2;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_A3;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_A4;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_A5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_A6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_AMUX;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_AO5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_AO6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_A_CY;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_A_XOR;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_B;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_B1;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_B2;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_B3;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_B4;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_B5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_B6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_BO5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_BO6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_B_CY;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_B_XOR;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_C;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_C1;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_C2;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_C3;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_C4;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_C5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_C6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_CLK;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_CO5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_CO6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_C_CY;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_C_XOR;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_D;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_D1;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_D2;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_D3;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_D4;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_D5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_D5Q;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_D6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_DMUX;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_DO5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_DO6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_DX;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_D_CY;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X0Y16_D_XOR;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_A;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_A1;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_A2;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_A3;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_A4;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_A5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_A6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_AO5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_AO6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_A_CY;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_A_XOR;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_B;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_B1;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_B2;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_B3;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_B4;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_B5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_B6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_BO5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_BO6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_B_CY;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_B_XOR;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_C;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_C1;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_C2;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_C3;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_C4;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_C5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_C6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_CO5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_CO6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_C_CY;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_C_XOR;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_D;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_D1;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_D2;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_D3;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_D4;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_D5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_D6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_DO5;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_DO6;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_D_CY;
  wire [0:0] CLBLL_L_X2Y16_SLICE_X1Y16_D_XOR;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_AO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_AO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A_XOR;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_BO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_BO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B_XOR;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_CO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_CO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C_XOR;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_DO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_DO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D_XOR;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_AMUX;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_AO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_AO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A_XOR;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_BO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_BO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B_XOR;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_CLK;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_CO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_CO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C_XOR;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D5Q;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_DMUX;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_DO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_DO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_DX;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D_XOR;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_A;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_A1;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_A2;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_A3;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_A4;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_A5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_A6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_AO5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_AO6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_A_CY;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_A_XOR;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_B;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_B1;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_B2;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_B3;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_B4;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_B5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_B6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_BO5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_BO6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_B_CY;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_B_XOR;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_C;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_C1;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_C2;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_C3;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_C4;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_C5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_C6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_CO5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_CO6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_C_CY;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_C_XOR;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_D;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_D1;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_D2;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_D3;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_D4;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_D5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_D6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_DO5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_DO6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_D_CY;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X0Y39_D_XOR;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_A;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_A1;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_A2;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_A3;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_A4;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_A5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_A6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_AMUX;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_AO5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_AO6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_A_CY;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_A_XOR;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_B;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_B1;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_B2;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_B3;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_B4;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_B5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_B6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_BO5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_BO6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_B_CY;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_B_XOR;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_C;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_C1;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_C2;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_C3;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_C4;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_C5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_C6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_CLK;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_CO5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_CO6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_C_CY;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_C_XOR;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_D;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_D1;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_D2;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_D3;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_D4;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_D5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_D5Q;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_D6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_DMUX;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_DO5;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_DO6;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_DX;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_D_CY;
  wire [0:0] CLBLL_L_X2Y39_SLICE_X1Y39_D_XOR;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_A;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_A1;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_A2;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_A3;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_A4;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_A5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_A6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_AMUX;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_AO5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_AO6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_A_CY;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_A_XOR;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_B;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_B1;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_B2;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_B3;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_B4;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_B5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_B6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_BMUX;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_BO5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_BO6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_B_CY;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_B_XOR;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_C;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_C1;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_C2;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_C3;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_C4;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_C5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_C6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_CO5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_CO6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_C_CY;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_C_XOR;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_D;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_D1;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_D2;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_D3;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_D4;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_D5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_D6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_DO5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_DO6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_D_CY;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X0Y5_D_XOR;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_A;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_A1;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_A2;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_A3;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_A4;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_A5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_A6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_AO5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_AO6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_A_CY;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_A_XOR;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_B;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_B1;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_B2;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_B3;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_B4;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_B5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_B6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_BO5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_BO6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_B_CY;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_B_XOR;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_C;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_C1;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_C2;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_C3;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_C4;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_C5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_C6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_CO5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_CO6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_C_CY;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_C_XOR;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_D;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_D1;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_D2;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_D3;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_D4;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_D5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_D6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_DO5;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_DO6;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_D_CY;
  wire [0:0] CLBLL_L_X2Y5_SLICE_X1Y5_D_XOR;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_A;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_A1;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_A2;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_A3;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_A4;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_A5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_A6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_AMUX;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_AO5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_AO6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_A_CY;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_A_XOR;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_B;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_B1;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_B2;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_B3;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_B4;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_B5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_B6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_BO5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_BO6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_B_CY;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_B_XOR;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_C;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_C1;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_C2;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_C3;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_C4;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_C5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_C6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_CLK;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_CO5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_CO6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_C_CY;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_C_XOR;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_D;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_D1;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_D2;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_D3;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_D4;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_D5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_D5Q;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_D6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_DMUX;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_DO5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_DO6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_DX;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_D_CY;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X0Y7_D_XOR;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_A;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_A1;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_A2;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_A3;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_A4;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_A5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_A6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_AO5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_AO6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_A_CY;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_A_XOR;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_B;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_B1;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_B2;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_B3;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_B4;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_B5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_B6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_BO5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_BO6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_B_CY;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_B_XOR;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_C;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_C1;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_C2;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_C3;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_C4;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_C5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_C6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_CO5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_CO6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_C_CY;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_C_XOR;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_D;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_D1;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_D2;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_D3;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_D4;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_D5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_D6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_DO5;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_DO6;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_D_CY;
  wire [0:0] CLBLL_L_X2Y7_SLICE_X1Y7_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_S1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_S1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S1;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBIN;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBOUT;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBOUTB;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBSTOPPED;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKIN1;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKIN2;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKINSEL;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKINSTOPPED;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT0;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT0B;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT1;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT1B;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT2;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT2B;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT3;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT3B;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR0;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR1;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR2;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR3;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR4;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR5;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR6;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DCLK;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DEN;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI0;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI1;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI10;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI11;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI12;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI13;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI14;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI15;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI2;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI3;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI4;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI5;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI6;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI7;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI8;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI9;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO0;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO1;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO10;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO11;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO12;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO13;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO14;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO15;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO2;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO3;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO4;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO5;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO6;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO7;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO8;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO9;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DRDY;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DWE;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_LOCKED;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSCLK;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSDONE;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSEN;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSINCDEC;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PWRDWN;
  wire [0:0] CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_RST;
  wire [0:0] LIOB33_SING_X0Y0_IOB_X0Y0_O;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y11_I;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y12_I;
  wire [0:0] LIOB33_X0Y17_IOB_X0Y18_O;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y19_O;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y20_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_O;
  wire [0:0] LIOB33_X0Y23_IOB_X0Y24_I;
  wire [0:0] LIOB33_X0Y25_IOB_X0Y25_I;
  wire [0:0] LIOB33_X0Y25_IOB_X0Y26_O;
  wire [0:0] LIOB33_X0Y27_IOB_X0Y28_O;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y3_O;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y4_O;
  wire [0:0] LIOB33_X0Y43_IOB_X0Y43_O;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y5_I;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y6_I;
  wire [0:0] LIOB33_X0Y7_IOB_X0Y7_I;
  wire [0:0] LIOB33_X0Y7_IOB_X0Y8_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y10_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y9_I;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_D1;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_OQ;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_T1;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_O;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_O;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_O;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_D1;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_OQ;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_T1;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_TQ;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y24_D;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y24_O;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y25_D;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y25_O;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y26_D1;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y26_OQ;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y26_T1;
  wire [0:0] LIOI3_X0Y25_OLOGIC_X0Y26_TQ;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_D1;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_OQ;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_T1;
  wire [0:0] LIOI3_X0Y27_OLOGIC_X0Y28_TQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_D1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_OQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_T1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_TQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_D1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_OQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_T1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_TQ;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y5_D;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y5_O;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_D;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_O;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_O;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y9_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y9_O;
  wire [0:0] RIOB33_X43Y25_IOB_X1Y26_I;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_D;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_O;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y5_SLICE_X0Y5_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y5_SLICE_X0Y5_DO5),
.O6(CLBLL_L_X2Y5_SLICE_X0Y5_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y5_SLICE_X0Y5_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y5_SLICE_X0Y5_CO5),
.O6(CLBLL_L_X2Y5_SLICE_X0Y5_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h00000f0f00330033)
  ) CLBLL_L_X2Y5_SLICE_X0Y5_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y11_IOB_X0Y11_I),
.I2(LIOB33_X0Y9_IOB_X0Y9_I),
.I3(LIOB33_X0Y11_IOB_X0Y12_I),
.I4(LIOB33_X0Y9_IOB_X0Y10_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y5_SLICE_X0Y5_BO5),
.O6(CLBLL_L_X2Y5_SLICE_X0Y5_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hfffffffdffffffff)
  ) CLBLL_L_X2Y5_SLICE_X0Y5_ALUT (
.I0(CLBLL_L_X2Y5_SLICE_X0Y5_BO6),
.I1(LIOB33_X0Y5_IOB_X0Y6_I),
.I2(LIOB33_X0Y5_IOB_X0Y5_I),
.I3(LIOB33_X0Y7_IOB_X0Y8_I),
.I4(LIOB33_X0Y7_IOB_X0Y7_I),
.I5(CLBLL_L_X2Y5_SLICE_X0Y5_BO5),
.O5(CLBLL_L_X2Y5_SLICE_X0Y5_AO5),
.O6(CLBLL_L_X2Y5_SLICE_X0Y5_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y5_SLICE_X1Y5_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y5_SLICE_X1Y5_DO5),
.O6(CLBLL_L_X2Y5_SLICE_X1Y5_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y5_SLICE_X1Y5_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y5_SLICE_X1Y5_CO5),
.O6(CLBLL_L_X2Y5_SLICE_X1Y5_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y5_SLICE_X1Y5_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y5_SLICE_X1Y5_BO5),
.O6(CLBLL_L_X2Y5_SLICE_X1Y5_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y5_SLICE_X1Y5_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y5_SLICE_X1Y5_AO5),
.O6(CLBLL_L_X2Y5_SLICE_X1Y5_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y7_SLICE_X0Y7_D5_FDRE (
.C(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.CE(1'b1),
.D(CLBLL_L_X2Y7_SLICE_X0Y7_AO5),
.Q(CLBLL_L_X2Y7_SLICE_X0Y7_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y7_SLICE_X0Y7_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y7_SLICE_X0Y7_DO5),
.O6(CLBLL_L_X2Y7_SLICE_X0Y7_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y7_SLICE_X0Y7_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y7_SLICE_X0Y7_CO5),
.O6(CLBLL_L_X2Y7_SLICE_X0Y7_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y7_SLICE_X0Y7_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y7_SLICE_X0Y7_BO5),
.O6(CLBLL_L_X2Y7_SLICE_X0Y7_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000f0f0f0f)
  ) CLBLL_L_X2Y7_SLICE_X0Y7_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y7_SLICE_X0Y7_D5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y7_SLICE_X0Y7_AO5),
.O6(CLBLL_L_X2Y7_SLICE_X0Y7_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y7_SLICE_X1Y7_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y7_SLICE_X1Y7_DO5),
.O6(CLBLL_L_X2Y7_SLICE_X1Y7_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y7_SLICE_X1Y7_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y7_SLICE_X1Y7_CO5),
.O6(CLBLL_L_X2Y7_SLICE_X1Y7_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y7_SLICE_X1Y7_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y7_SLICE_X1Y7_BO5),
.O6(CLBLL_L_X2Y7_SLICE_X1Y7_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y7_SLICE_X1Y7_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y7_SLICE_X1Y7_AO5),
.O6(CLBLL_L_X2Y7_SLICE_X1Y7_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y16_SLICE_X0Y16_D5_FDRE (
.C(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_O),
.CE(1'b1),
.D(CLBLL_L_X2Y16_SLICE_X0Y16_AO5),
.Q(CLBLL_L_X2Y16_SLICE_X0Y16_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y16_SLICE_X0Y16_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y16_SLICE_X0Y16_DO5),
.O6(CLBLL_L_X2Y16_SLICE_X0Y16_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y16_SLICE_X0Y16_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y16_SLICE_X0Y16_CO5),
.O6(CLBLL_L_X2Y16_SLICE_X0Y16_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y16_SLICE_X0Y16_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y16_SLICE_X0Y16_BO5),
.O6(CLBLL_L_X2Y16_SLICE_X0Y16_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000f0f0f0f)
  ) CLBLL_L_X2Y16_SLICE_X0Y16_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y16_SLICE_X0Y16_D5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y16_SLICE_X0Y16_AO5),
.O6(CLBLL_L_X2Y16_SLICE_X0Y16_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y16_SLICE_X1Y16_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y16_SLICE_X1Y16_DO5),
.O6(CLBLL_L_X2Y16_SLICE_X1Y16_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y16_SLICE_X1Y16_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y16_SLICE_X1Y16_CO5),
.O6(CLBLL_L_X2Y16_SLICE_X1Y16_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y16_SLICE_X1Y16_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y16_SLICE_X1Y16_BO5),
.O6(CLBLL_L_X2Y16_SLICE_X1Y16_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y16_SLICE_X1Y16_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y16_SLICE_X1Y16_AO5),
.O6(CLBLL_L_X2Y16_SLICE_X1Y16_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y23_SLICE_X0Y23_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X0Y23_DO5),
.O6(CLBLL_L_X2Y23_SLICE_X0Y23_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y23_SLICE_X0Y23_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X0Y23_CO5),
.O6(CLBLL_L_X2Y23_SLICE_X0Y23_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y23_SLICE_X0Y23_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X0Y23_BO5),
.O6(CLBLL_L_X2Y23_SLICE_X0Y23_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y23_SLICE_X0Y23_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X0Y23_AO5),
.O6(CLBLL_L_X2Y23_SLICE_X0Y23_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y23_SLICE_X1Y23_D5_FDRE (
.C(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_O),
.CE(1'b1),
.D(CLBLL_L_X2Y23_SLICE_X1Y23_AO5),
.Q(CLBLL_L_X2Y23_SLICE_X1Y23_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y23_SLICE_X1Y23_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X1Y23_DO5),
.O6(CLBLL_L_X2Y23_SLICE_X1Y23_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y23_SLICE_X1Y23_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X1Y23_CO5),
.O6(CLBLL_L_X2Y23_SLICE_X1Y23_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y23_SLICE_X1Y23_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X1Y23_BO5),
.O6(CLBLL_L_X2Y23_SLICE_X1Y23_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000f0f0f0f)
  ) CLBLL_L_X2Y23_SLICE_X1Y23_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y23_SLICE_X1Y23_D5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X1Y23_AO5),
.O6(CLBLL_L_X2Y23_SLICE_X1Y23_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y39_SLICE_X0Y39_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y39_SLICE_X0Y39_DO5),
.O6(CLBLL_L_X2Y39_SLICE_X0Y39_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y39_SLICE_X0Y39_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y39_SLICE_X0Y39_CO5),
.O6(CLBLL_L_X2Y39_SLICE_X0Y39_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y39_SLICE_X0Y39_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y39_SLICE_X0Y39_BO5),
.O6(CLBLL_L_X2Y39_SLICE_X0Y39_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y39_SLICE_X0Y39_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y39_SLICE_X0Y39_AO5),
.O6(CLBLL_L_X2Y39_SLICE_X0Y39_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D5FF" *)
  FDRE #(
    .INIT(1),
    .IS_C_INVERTED(0)
  ) CLBLL_L_X2Y39_SLICE_X1Y39_D5_FDRE (
.C(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O),
.CE(1'b1),
.D(CLBLL_L_X2Y39_SLICE_X1Y39_AO5),
.Q(CLBLL_L_X2Y39_SLICE_X1Y39_D5Q),
.R(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y39_SLICE_X1Y39_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y39_SLICE_X1Y39_DO5),
.O6(CLBLL_L_X2Y39_SLICE_X1Y39_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y39_SLICE_X1Y39_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y39_SLICE_X1Y39_CO5),
.O6(CLBLL_L_X2Y39_SLICE_X1Y39_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y39_SLICE_X1Y39_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y39_SLICE_X1Y39_BO5),
.O6(CLBLL_L_X2Y39_SLICE_X1Y39_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h000000000f0f0f0f)
  ) CLBLL_L_X2Y39_SLICE_X1Y39_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(CLBLL_L_X2Y39_SLICE_X1Y39_D5Q),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y39_SLICE_X1Y39_AO5),
.O6(CLBLL_L_X2Y39_SLICE_X1Y39_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT0),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT1),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT2),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT3),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "MMCME2_ADV" *)
  MMCME2_ADV #(
    .BANDWIDTH("OPTIMIZED"),
    .CLKFBOUT_MULT_F(10.500),
    .CLKFBOUT_PHASE(0.000),
    .CLKIN1_PERIOD(11.667),
    .CLKIN2_PERIOD(11.667),
    .CLKOUT0_DIVIDE_F(12.500),
    .CLKOUT0_DUTY_CYCLE(0.500),
    .CLKOUT0_PHASE(43.200),
    .CLKOUT1_DIVIDE(32),
    .CLKOUT1_DUTY_CYCLE(0.5312),
    .CLKOUT1_PHASE(90.000),
    .CLKOUT2_DIVIDE(48),
    .CLKOUT2_DUTY_CYCLE(0.5000),
    .CLKOUT2_PHASE(135.000),
    .CLKOUT3_DIVIDE(64),
    .CLKOUT3_DUTY_CYCLE(0.5000),
    .CLKOUT3_PHASE(45.000),
    .CLKOUT4_DIVIDE(1),
    .CLKOUT4_DUTY_CYCLE(0.500),
    .CLKOUT4_PHASE(0.000),
    .CLKOUT5_DIVIDE(1),
    .CLKOUT5_DUTY_CYCLE(0.500),
    .CLKOUT5_PHASE(0.000),
    .CLKOUT6_DIVIDE(1),
    .CLKOUT6_DUTY_CYCLE(0.500),
    .CLKOUT6_PHASE(0.000),
    .COMPENSATION("INTERNAL"),
    .DIVCLK_DIVIDE(1),
    .IS_CLKINSEL_INVERTED(1'b1),
    .IS_PSEN_INVERTED(1'b1),
    .IS_PSINCDEC_INVERTED(1'b1),
    .IS_PWRDWN_INVERTED(1'b1),
    .IS_RST_INVERTED(1'b0),
    .SS_EN("FALSE"),
    .SS_MODE("CENTER_HIGH"),
    .SS_MOD_PERIOD(10000),
    .STARTUP_WAIT("FALSE")
  ) CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_MMCME2_ADV (
.CLKFBIN(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBOUT),
.CLKFBOUT(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBOUT),
.CLKFBOUTB(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBOUTB),
.CLKFBSTOPPED(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBSTOPPED),
.CLKIN1(RIOB33_X43Y25_IOB_X1Y26_I),
.CLKIN2(RIOB33_X43Y25_IOB_X1Y26_I),
.CLKINSEL(1'b1),
.CLKINSTOPPED(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKINSTOPPED),
.CLKOUT0(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT0),
.CLKOUT0B(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT0B),
.CLKOUT1(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT1),
.CLKOUT1B(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT1B),
.CLKOUT2(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT2),
.CLKOUT2B(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT2B),
.CLKOUT3(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT3),
.CLKOUT3B(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT3B),
.DADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.DCLK(1'b0),
.DEN(1'b0),
.DI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.DO({CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO15, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO14, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO13, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO12, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO11, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO10, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO9, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO8, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO7, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO6, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO5, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO4, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO3, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO2, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO1, CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DO0}),
.DRDY(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DRDY),
.DWE(1'b0),
.LOCKED(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_LOCKED),
.PSCLK(1'b0),
.PSDONE(CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSDONE),
.PSEN(1'b1),
.PSINCDEC(1'b1),
.PWRDWN(1'b1),
.RST(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y1_OBUF (
.I(CLBLL_L_X2Y5_SLICE_X0Y5_AO6),
.O(led[7])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y3_IOB_X0Y3_OBUF (
.I(CLBLL_L_X2Y7_SLICE_X0Y7_D5Q),
.O(led[0])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y3_IOB_X0Y4_OBUF (
.I(1'b0),
.O(led[5])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y5_IOB_X0Y5_IBUF (
.I(sw[6]),
.O(LIOB33_X0Y5_IOB_X0Y5_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y5_IOB_X0Y6_IBUF (
.I(sw[7]),
.O(LIOB33_X0Y5_IOB_X0Y6_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y7_IOB_X0Y7_IBUF (
.I(sw[4]),
.O(LIOB33_X0Y7_IOB_X0Y7_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y7_IOB_X0Y8_IBUF (
.I(sw[5]),
.O(LIOB33_X0Y7_IOB_X0Y8_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y9_IOB_X0Y9_IBUF (
.I(sw[3]),
.O(LIOB33_X0Y9_IOB_X0Y9_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y9_IOB_X0Y10_IBUF (
.I(sw[2]),
.O(LIOB33_X0Y9_IOB_X0Y10_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y11_IOB_X0Y11_IBUF (
.I(sw[0]),
.O(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y11_IOB_X0Y12_IBUF (
.I(sw[1]),
.O(LIOB33_X0Y11_IOB_X0Y12_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y17_IOB_X0Y18_OBUF (
.I(1'b0),
.O(led[4])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y19_IOB_X0Y19_OBUF (
.I(CLBLL_L_X2Y23_SLICE_X1Y23_D5Q),
.O(led[3])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y19_IOB_X0Y20_OBUF (
.I(CLBLL_L_X2Y16_SLICE_X0Y16_D5Q),
.O(led[2])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y23_IOB_X0Y24_IBUF (
.I(jc3),
.O(LIOB33_X0Y23_IOB_X0Y24_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y25_IOB_X0Y25_IBUF (
.I(jc1),
.O(LIOB33_X0Y25_IOB_X0Y25_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y25_IOB_X0Y26_OBUF (
.I(LIOB33_X0Y23_IOB_X0Y24_I),
.O(jc4)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y27_IOB_X0Y28_OBUF (
.I(LIOB33_X0Y25_IOB_X0Y25_I),
.O(jc2)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y43_IOB_X0Y43_OBUF (
.I(CLBLL_L_X2Y39_SLICE_X1Y39_D5Q),
.O(led[1])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y0_IOB_X0Y0_OBUF (
.I(1'b0),
.O(led[6])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y25_IOB_X1Y26_IBUF (
.I(clk),
.O(RIOB33_X43Y25_IOB_X1Y26_I)
  );
  assign CLBLL_L_X2Y5_SLICE_X0Y5_COUT = CLBLL_L_X2Y5_SLICE_X0Y5_D_CY;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_A = CLBLL_L_X2Y5_SLICE_X0Y5_AO6;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_B = CLBLL_L_X2Y5_SLICE_X0Y5_BO6;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_C = CLBLL_L_X2Y5_SLICE_X0Y5_CO6;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_D = CLBLL_L_X2Y5_SLICE_X0Y5_DO6;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_AMUX = CLBLL_L_X2Y5_SLICE_X0Y5_AO6;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_BMUX = CLBLL_L_X2Y5_SLICE_X0Y5_BO5;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_COUT = CLBLL_L_X2Y5_SLICE_X1Y5_D_CY;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_A = CLBLL_L_X2Y5_SLICE_X1Y5_AO6;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_B = CLBLL_L_X2Y5_SLICE_X1Y5_BO6;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_C = CLBLL_L_X2Y5_SLICE_X1Y5_CO6;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_D = CLBLL_L_X2Y5_SLICE_X1Y5_DO6;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_COUT = CLBLL_L_X2Y7_SLICE_X0Y7_D_CY;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_A = CLBLL_L_X2Y7_SLICE_X0Y7_AO6;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_B = CLBLL_L_X2Y7_SLICE_X0Y7_BO6;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_C = CLBLL_L_X2Y7_SLICE_X0Y7_CO6;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_D = CLBLL_L_X2Y7_SLICE_X0Y7_DO6;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_AMUX = CLBLL_L_X2Y7_SLICE_X0Y7_AO5;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_DMUX = CLBLL_L_X2Y7_SLICE_X0Y7_D5Q;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_COUT = CLBLL_L_X2Y7_SLICE_X1Y7_D_CY;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_A = CLBLL_L_X2Y7_SLICE_X1Y7_AO6;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_B = CLBLL_L_X2Y7_SLICE_X1Y7_BO6;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_C = CLBLL_L_X2Y7_SLICE_X1Y7_CO6;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_D = CLBLL_L_X2Y7_SLICE_X1Y7_DO6;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_COUT = CLBLL_L_X2Y16_SLICE_X0Y16_D_CY;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_A = CLBLL_L_X2Y16_SLICE_X0Y16_AO6;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_B = CLBLL_L_X2Y16_SLICE_X0Y16_BO6;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_C = CLBLL_L_X2Y16_SLICE_X0Y16_CO6;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_D = CLBLL_L_X2Y16_SLICE_X0Y16_DO6;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_AMUX = CLBLL_L_X2Y16_SLICE_X0Y16_AO5;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_DMUX = CLBLL_L_X2Y16_SLICE_X0Y16_D5Q;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_COUT = CLBLL_L_X2Y16_SLICE_X1Y16_D_CY;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_A = CLBLL_L_X2Y16_SLICE_X1Y16_AO6;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_B = CLBLL_L_X2Y16_SLICE_X1Y16_BO6;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_C = CLBLL_L_X2Y16_SLICE_X1Y16_CO6;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_D = CLBLL_L_X2Y16_SLICE_X1Y16_DO6;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_COUT = CLBLL_L_X2Y23_SLICE_X0Y23_D_CY;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_A = CLBLL_L_X2Y23_SLICE_X0Y23_AO6;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_B = CLBLL_L_X2Y23_SLICE_X0Y23_BO6;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_C = CLBLL_L_X2Y23_SLICE_X0Y23_CO6;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_D = CLBLL_L_X2Y23_SLICE_X0Y23_DO6;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_COUT = CLBLL_L_X2Y23_SLICE_X1Y23_D_CY;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_A = CLBLL_L_X2Y23_SLICE_X1Y23_AO6;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_B = CLBLL_L_X2Y23_SLICE_X1Y23_BO6;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_C = CLBLL_L_X2Y23_SLICE_X1Y23_CO6;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_D = CLBLL_L_X2Y23_SLICE_X1Y23_DO6;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_AMUX = CLBLL_L_X2Y23_SLICE_X1Y23_AO5;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_DMUX = CLBLL_L_X2Y23_SLICE_X1Y23_D5Q;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_COUT = CLBLL_L_X2Y39_SLICE_X0Y39_D_CY;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_A = CLBLL_L_X2Y39_SLICE_X0Y39_AO6;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_B = CLBLL_L_X2Y39_SLICE_X0Y39_BO6;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_C = CLBLL_L_X2Y39_SLICE_X0Y39_CO6;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_D = CLBLL_L_X2Y39_SLICE_X0Y39_DO6;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_COUT = CLBLL_L_X2Y39_SLICE_X1Y39_D_CY;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_A = CLBLL_L_X2Y39_SLICE_X1Y39_AO6;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_B = CLBLL_L_X2Y39_SLICE_X1Y39_BO6;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_C = CLBLL_L_X2Y39_SLICE_X1Y39_CO6;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_D = CLBLL_L_X2Y39_SLICE_X1Y39_DO6;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_AMUX = CLBLL_L_X2Y39_SLICE_X1Y39_AO5;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_DMUX = CLBLL_L_X2Y39_SLICE_X1Y39_D5Q;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_OQ = CLBLL_L_X2Y5_SLICE_X0Y5_AO6;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_TQ = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_OQ = 1'b0;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_TQ = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_OQ = CLBLL_L_X2Y7_SLICE_X0Y7_D5Q;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_TQ = 1'b1;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_O = LIOB33_X0Y5_IOB_X0Y6_I;
  assign LIOI3_X0Y5_ILOGIC_X0Y5_O = LIOB33_X0Y5_IOB_X0Y5_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_O = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y9_O = LIOB33_X0Y9_IOB_X0Y9_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_O = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_O = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_OQ = 1'b0;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_TQ = 1'b1;
  assign LIOI3_X0Y23_ILOGIC_X0Y24_O = LIOB33_X0Y23_IOB_X0Y24_I;
  assign LIOI3_X0Y25_ILOGIC_X0Y25_O = LIOB33_X0Y25_IOB_X0Y25_I;
  assign LIOI3_X0Y25_OLOGIC_X0Y26_OQ = LIOB33_X0Y23_IOB_X0Y24_I;
  assign LIOI3_X0Y25_OLOGIC_X0Y26_TQ = 1'b1;
  assign LIOI3_X0Y27_OLOGIC_X0Y28_OQ = LIOB33_X0Y25_IOB_X0Y25_I;
  assign LIOI3_X0Y27_OLOGIC_X0Y28_TQ = 1'b1;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_OQ = 1'b0;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_O = LIOB33_X0Y7_IOB_X0Y8_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_O = LIOB33_X0Y7_IOB_X0Y7_I;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_OQ = CLBLL_L_X2Y16_SLICE_X0Y16_D5Q;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_OQ = CLBLL_L_X2Y23_SLICE_X1Y23_D5Q;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ = CLBLL_L_X2Y39_SLICE_X1Y39_D5Q;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ = 1'b1;
  assign RIOI3_X43Y25_ILOGIC_X1Y26_O = RIOB33_X43Y25_IOB_X1Y26_I;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_D1 = CLBLL_L_X2Y16_SLICE_X0Y16_D5Q;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_T1 = 1'b1;
  assign LIOB33_X0Y1_IOB_X0Y1_O = CLBLL_L_X2Y5_SLICE_X0Y5_AO6;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_D = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y9_D = LIOB33_X0Y9_IOB_X0Y9_I;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_A1 = CLBLL_L_X2Y5_SLICE_X0Y5_BO6;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_A2 = LIOB33_X0Y5_IOB_X0Y6_I;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_A3 = LIOB33_X0Y5_IOB_X0Y5_I;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_A4 = LIOB33_X0Y7_IOB_X0Y8_I;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_A5 = LIOB33_X0Y7_IOB_X0Y7_I;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_A6 = CLBLL_L_X2Y5_SLICE_X0Y5_BO5;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_B1 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_B2 = LIOB33_X0Y11_IOB_X0Y11_I;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_B3 = LIOB33_X0Y9_IOB_X0Y9_I;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_B4 = LIOB33_X0Y11_IOB_X0Y12_I;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_B5 = LIOB33_X0Y9_IOB_X0Y10_I;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_B6 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI2 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI3 = 1'b0;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_C1 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_C2 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_C3 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_C4 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_C5 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_C6 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI4 = 1'b0;
  assign LIOB33_SING_X0Y0_IOB_X0Y0_O = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI5 = 1'b0;
  assign LIOI3_X0Y25_OLOGIC_X0Y26_D1 = LIOB33_X0Y23_IOB_X0Y24_I;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI6 = 1'b0;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_D1 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_D2 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_D3 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_D4 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_D5 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X0Y5_D6 = 1'b1;
  assign LIOI3_X0Y25_OLOGIC_X0Y26_T1 = 1'b1;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_D1 = 1'b0;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_T1 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_A1 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_A2 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_A3 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_A4 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_A5 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_A6 = 1'b1;
  assign LIOB33_X0Y17_IOB_X0Y18_O = 1'b0;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_B1 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_B2 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_B3 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_B4 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_B5 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_B6 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_C1 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_C2 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_C3 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_C4 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_C5 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_C6 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_D1 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_D2 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_D3 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_D4 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_D5 = 1'b1;
  assign CLBLL_L_X2Y5_SLICE_X1Y5_D6 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S1 = 1'b1;
  assign LIOB33_X0Y3_IOB_X0Y3_O = CLBLL_L_X2Y7_SLICE_X0Y7_D5Q;
  assign LIOB33_X0Y3_IOB_X0Y4_O = 1'b0;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_D = LIOB33_X0Y5_IOB_X0Y6_I;
  assign LIOI3_X0Y5_ILOGIC_X0Y5_D = LIOB33_X0Y5_IOB_X0Y5_I;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_D1 = CLBLL_L_X2Y23_SLICE_X1Y23_D5Q;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_T1 = 1'b1;
  assign LIOB33_X0Y25_IOB_X0Y26_O = LIOB33_X0Y23_IOB_X0Y24_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_S1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_S1 = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_D1 = 1'b0;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_D = LIOB33_X0Y7_IOB_X0Y7_I;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_T1 = 1'b1;
  assign LIOI3_X0Y25_ILOGIC_X0Y25_D = LIOB33_X0Y25_IOB_X0Y25_I;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_D1 = CLBLL_L_X2Y7_SLICE_X0Y7_D5Q;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_T1 = 1'b1;
  assign RIOI3_X43Y25_ILOGIC_X1Y26_D = RIOB33_X43Y25_IOB_X1Y26_I;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1 = CLBLL_L_X2Y39_SLICE_X1Y39_D5Q;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_A1 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_A2 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_A3 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_A4 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_A5 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_A6 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_B1 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_B2 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_B3 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_B4 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_B5 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_B6 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_C1 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_C2 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_C3 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_C4 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_C5 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_C6 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_D1 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_D2 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_D3 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_A1 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_A2 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_D6 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_A3 = CLBLL_L_X2Y16_SLICE_X0Y16_D5Q;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_A4 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_A5 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_A6 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_D4 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X0Y39_D5 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_B1 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_B2 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_B4 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_B5 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_B6 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_B3 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_C1 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_C2 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_C3 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_C4 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_C5 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_C6 = 1'b1;
  assign LIOB33_X0Y19_IOB_X0Y19_O = CLBLL_L_X2Y23_SLICE_X1Y23_D5Q;
  assign LIOB33_X0Y19_IOB_X0Y20_O = CLBLL_L_X2Y16_SLICE_X0Y16_D5Q;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_A1 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_A2 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_D1 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_D2 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_D3 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_D4 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_D5 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_D6 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_A3 = CLBLL_L_X2Y39_SLICE_X1Y39_D5Q;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_A4 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_DX = CLBLL_L_X2Y16_SLICE_X0Y16_AO5;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_A5 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_A6 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_B1 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_B2 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_B3 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_B4 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_B5 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_B6 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_C1 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_C2 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_C3 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_C4 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_C5 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_C6 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_D1 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_D2 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_D3 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_A1 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_A2 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_A3 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_A4 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_A5 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_DX = CLBLL_L_X2Y39_SLICE_X1Y39_AO5;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_A6 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_D4 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_D5 = 1'b1;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_D6 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_B1 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_B2 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_B3 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_B4 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_B5 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_B6 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_C1 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_C2 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_C3 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_C4 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_C5 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_C6 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_D1 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_D2 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_D3 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_D4 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_D5 = 1'b1;
  assign CLBLL_L_X2Y16_SLICE_X1Y16_D6 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_A1 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_A2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_A3 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_A4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_A5 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_A6 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_B1 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_B2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_B3 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_B4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_B5 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_B6 = 1'b1;
  assign LIOB33_X0Y27_IOB_X0Y28_O = LIOB33_X0Y25_IOB_X0Y25_I;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_C1 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_C2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_C3 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_C4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_C5 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_C6 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_D1 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_D2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_D3 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_D4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_D5 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_D6 = 1'b1;
  assign LIOI3_X0Y23_ILOGIC_X0Y24_D = LIOB33_X0Y23_IOB_X0Y24_I;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_D1 = CLBLL_L_X2Y5_SLICE_X0Y5_AO6;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_T1 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_A1 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_A2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_A3 = CLBLL_L_X2Y23_SLICE_X1Y23_D5Q;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_A4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_A5 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_A6 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_B1 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_B2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_B3 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_B4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_B5 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_B6 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_C1 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_C2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_C3 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_C4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_C5 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_C6 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_D1 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_D2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_D3 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_D4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_D5 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_D6 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_DX = CLBLL_L_X2Y23_SLICE_X1Y23_AO5;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_D = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_D = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_D = LIOB33_X0Y7_IOB_X0Y8_I;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_A1 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_A2 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_A3 = CLBLL_L_X2Y7_SLICE_X0Y7_D5Q;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_A4 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_A5 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_A6 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_B1 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_B2 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_B3 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_B4 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_B5 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_B6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_C1 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_C2 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_C3 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_C4 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_C5 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_C6 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_D1 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_D2 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_D3 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_D4 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_D5 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_D6 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_DX = CLBLL_L_X2Y7_SLICE_X0Y7_AO5;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_A1 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_A2 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_A3 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_A4 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_A5 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_A6 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBIN = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKFBOUT;
  assign LIOB33_X0Y43_IOB_X0Y43_O = CLBLL_L_X2Y39_SLICE_X1Y39_D5Q;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_B1 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_B2 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_B3 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_B4 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_B5 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_B6 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKIN1 = RIOB33_X43Y25_IOB_X1Y26_I;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKIN2 = RIOB33_X43Y25_IOB_X1Y26_I;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKINSEL = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_C1 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_C2 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_C3 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_C4 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_C5 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_C6 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR0 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR1 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR2 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR3 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR4 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR5 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DADDR6 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DCLK = 1'b0;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_D1 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_D2 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_D3 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_D4 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_D5 = 1'b1;
  assign CLBLL_L_X2Y7_SLICE_X1Y7_D6 = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DEN = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI0 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI1 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI11 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI12 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI13 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI14 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI15 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI7 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI8 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI9 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DI10 = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_DWE = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSCLK = 1'b0;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSEN = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PSINCDEC = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_PWRDWN = 1'b1;
  assign CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_RST = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOI3_X0Y27_OLOGIC_X0Y28_D1 = LIOB33_X0Y25_IOB_X0Y25_I;
  assign LIOI3_X0Y27_OLOGIC_X0Y28_T1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0 = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT0;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I0 = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_I0 = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT2;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_I1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_I0 = CMT_TOP_L_LOWER_B_X106Y9_MMCME2_ADV_X1Y0_CLKOUT3;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_I1 = 1'b1;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_D1 = 1'b0;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_CLK = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y11_O;
  assign CLBLL_L_X2Y39_SLICE_X1Y39_CLK = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O;
  assign CLBLL_L_X2Y16_SLICE_X0Y16_CLK = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y10_O;
  assign CLBLL_L_X2Y7_SLICE_X0Y7_CLK = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
endmodule
