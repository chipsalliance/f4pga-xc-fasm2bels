module top(
  input LIOB33_SING_X0Y0_IOB_X0Y0_IPAD,
  input LIOB33_X0Y1_IOB_X0Y1_IPAD,
  output LIOB33_X0Y1_IOB_X0Y2_OPAD
  );
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_A;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_A1;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_A2;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_A3;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_A4;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_A5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_A6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_AO5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_AO6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_A_CY;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_A_XOR;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_B;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_B1;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_B2;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_B3;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_B4;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_B5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_B6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_BO5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_BO6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_B_CY;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_B_XOR;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_C;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_C1;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_C2;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_C3;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_C4;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_C5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_C6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_CO5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_CO6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_C_CY;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_C_XOR;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_D;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_D1;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_D2;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_D3;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_D4;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_D5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_D6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_DO5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_DO6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_D_CY;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X0Y1_D_XOR;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_A;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_A1;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_A2;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_A3;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_A4;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_A5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_A6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_AO5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_AO6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_A_CY;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_A_XOR;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_B;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_B1;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_B2;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_B3;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_B4;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_B5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_B6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_BO5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_BO6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_B_CY;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_B_XOR;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_C;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_C1;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_C2;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_C3;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_C4;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_C5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_C6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_CO5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_CO6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_C_CY;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_C_XOR;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_D;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_D1;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_D2;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_D3;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_D4;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_D5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_D6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_DO5;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_DO6;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_D_CY;
  wire [0:0] CLBLL_L_X2Y1_SLICE_X1Y1_D_XOR;
  wire [0:0] LIOB33_SING_X0Y0_IOB_X0Y0_I;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_I;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y2_O;
  wire [0:0] LIOI3_SING_X0Y0_ILOGIC_X0Y0_D;
  wire [0:0] LIOI3_SING_X0Y0_ILOGIC_X0Y0_O;
  wire [0:0] LIOI3_X0Y1_ILOGIC_X0Y1_D;
  wire [0:0] LIOI3_X0Y1_ILOGIC_X0Y1_O;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_TQ;


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y1_SLICE_X0Y1_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y1_SLICE_X0Y1_DO5),
.O6(CLBLL_L_X2Y1_SLICE_X0Y1_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y1_SLICE_X0Y1_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y1_SLICE_X0Y1_CO5),
.O6(CLBLL_L_X2Y1_SLICE_X0Y1_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y1_SLICE_X0Y1_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y1_SLICE_X0Y1_BO5),
.O6(CLBLL_L_X2Y1_SLICE_X0Y1_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'hf0f00000f0f00000)
  ) CLBLL_L_X2Y1_SLICE_X0Y1_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y1_IOB_X0Y1_I),
.I3(1'b1),
.I4(LIOB33_SING_X0Y0_IOB_X0Y0_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y1_SLICE_X0Y1_AO5),
.O6(CLBLL_L_X2Y1_SLICE_X0Y1_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y1_SLICE_X1Y1_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y1_SLICE_X1Y1_DO5),
.O6(CLBLL_L_X2Y1_SLICE_X1Y1_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y1_SLICE_X1Y1_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y1_SLICE_X1Y1_CO5),
.O6(CLBLL_L_X2Y1_SLICE_X1Y1_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y1_SLICE_X1Y1_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y1_SLICE_X1Y1_BO5),
.O6(CLBLL_L_X2Y1_SLICE_X1Y1_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y1_SLICE_X1Y1_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y1_SLICE_X1Y1_AO5),
.O6(CLBLL_L_X2Y1_SLICE_X1Y1_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y1_IOB_X0Y1_IBUF (
.I(LIOB33_X0Y1_IOB_X0Y1_IPAD),
.O(LIOB33_X0Y1_IOB_X0Y1_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y2_OBUF (
.I(CLBLL_L_X2Y1_SLICE_X0Y1_AO6),
.O(LIOB33_X0Y1_IOB_X0Y2_OPAD)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_SING_X0Y0_IOB_X0Y0_IBUF (
.I(LIOB33_SING_X0Y0_IOB_X0Y0_IPAD),
.O(LIOB33_SING_X0Y0_IOB_X0Y0_I)
  );
  assign CLBLL_L_X2Y1_SLICE_X0Y1_A = CLBLL_L_X2Y1_SLICE_X0Y1_AO6;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_B = CLBLL_L_X2Y1_SLICE_X0Y1_BO6;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_C = CLBLL_L_X2Y1_SLICE_X0Y1_CO6;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_D = CLBLL_L_X2Y1_SLICE_X0Y1_DO6;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_A = CLBLL_L_X2Y1_SLICE_X1Y1_AO6;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_B = CLBLL_L_X2Y1_SLICE_X1Y1_BO6;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_C = CLBLL_L_X2Y1_SLICE_X1Y1_CO6;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_D = CLBLL_L_X2Y1_SLICE_X1Y1_DO6;
  assign LIOI3_X0Y1_ILOGIC_X0Y1_O = LIOB33_X0Y1_IOB_X0Y1_I;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_OQ = CLBLL_L_X2Y1_SLICE_X0Y1_AO6;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_TQ = 1'b1;
  assign LIOI3_SING_X0Y0_ILOGIC_X0Y0_O = LIOB33_SING_X0Y0_IOB_X0Y0_I;
  assign LIOB33_X0Y1_IOB_X0Y2_O = CLBLL_L_X2Y1_SLICE_X0Y1_AO6;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_D1 = CLBLL_L_X2Y1_SLICE_X0Y1_AO6;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_A1 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_A2 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_A3 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_A4 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_A5 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_A6 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_B1 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_B2 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_B3 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_B4 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_B5 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_B6 = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_T1 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_C1 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_C2 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_C3 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_C4 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_C5 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_C6 = 1'b1;
  assign LIOI3_SING_X0Y0_ILOGIC_X0Y0_D = LIOB33_SING_X0Y0_IOB_X0Y0_I;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_D1 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_D2 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_D3 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_D4 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_D5 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X1Y1_D6 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_A1 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_A2 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_A3 = LIOB33_X0Y1_IOB_X0Y1_I;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_A4 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_A5 = LIOB33_SING_X0Y0_IOB_X0Y0_I;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_A6 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_B1 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_B2 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_B3 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_B4 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_B5 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_B6 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_C1 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_C2 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_C3 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_C4 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_C5 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_C6 = 1'b1;
  assign LIOI3_X0Y1_ILOGIC_X0Y1_D = LIOB33_X0Y1_IOB_X0Y1_I;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_D1 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_D2 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_D3 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_D4 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_D5 = 1'b1;
  assign CLBLL_L_X2Y1_SLICE_X0Y1_D6 = 1'b1;
endmodule

