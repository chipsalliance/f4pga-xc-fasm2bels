// Copyright (C) 2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC

module top(
  input GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_IPAD_RX_N,
  input GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_IPAD_RX_P,
  input GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y0_IPAD_N,
  input GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y0_IPAD_P,
  input GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y1_IPAD_N,
  input GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y1_IPAD_P,
  input test_in,
  output GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_OPAD_TX_N,
  output GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_OPAD_TX_P,
  output test_out
  );
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_CFGRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_CLKRSVD0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_CLKRSVD1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONFIFORESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITORCLK;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT10;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT11;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT12;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT13;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT14;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT5;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT6;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT7;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT8;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT9;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR5;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR6;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR7;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR8;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPCLK;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI10;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI11;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI12;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI13;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI14;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI15;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI5;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI6;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI7;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI8;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI9;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO10;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO11;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO12;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO13;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO14;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO15;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO5;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO6;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO7;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO8;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO9;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPRDY;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPWE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_EYESCANDATAERROR;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_EYESCANMODE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_EYESCANRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_EYESCANTRIGGER;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRESETSEL;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD10;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD11;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD12;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD13;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD14;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD15;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD5;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD6;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD7;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD8;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD9;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRXRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTTXRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_LOOPBACK0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_LOOPBACK1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_LOOPBACK2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN10;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN11;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN12;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN13;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN14;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN15;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN5;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN6;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN7;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN8;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN9;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT10;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT11;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT12;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT13;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT14;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT15;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT5;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT6;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT7;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT8;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT9;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PHYSTATUS;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PMARSVDIN0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PMARSVDIN1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PMARSVDIN2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PMARSVDIN3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PMARSVDIN4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PMARSVDOUT0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PMARSVDOUT1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RESETOVRD;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RX8B10BEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST10;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST11;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST12;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST13;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST5;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST6;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST7;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST8;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST9;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXBUFRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXBUFSTATUS0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXBUFSTATUS1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXBUFSTATUS2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXBYTEISALIGNED;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXBYTEREALIGN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCDRFREQRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCDRHOLD;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCDRLOCK;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCDROVRDEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCDRRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCDRRESETRSV;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHANBONDSEQ;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHANISALIGNED;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHANREALIGN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISCOMMA0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISCOMMA1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISCOMMA2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISCOMMA3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISK0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISK1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISK2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISK3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDI0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDI1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDI2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDI3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDLEVEL0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDLEVEL1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDLEVEL2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDMASTER;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDO0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDO1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDO2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDO3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDSLAVE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCLKCORCNT0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCLKCORCNT1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCOMINITDET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCOMMADET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCOMMADETEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCOMSASDET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCOMWAKEDET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA10;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA11;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA12;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA13;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA14;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA15;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA16;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA17;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA18;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA19;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA20;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA21;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA22;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA23;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA24;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA25;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA26;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA27;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA28;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA29;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA30;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA31;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA5;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA6;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA7;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA8;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA9;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATAVALID0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATAVALID1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDDIEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDFEXYDEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDISPERR0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDISPERR1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDISPERR2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDISPERR3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDLYBYPASS;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDLYEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDLYOVRDEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDLYSRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDLYSRESETDONE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXELECIDLE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXELECIDLEMODE0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXELECIDLEMODE1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXGEARBOXSLIP;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXHEADER0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXHEADER1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXHEADER2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXHEADERVALID;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXLPMHFHOLD;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXLPMHFOVRDEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXLPMLFHOLD;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXLPMLFOVRDEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXLPMOSINTNTRLEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXLPMRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXMCOMMAALIGNEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXNOTINTABLE0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXNOTINTABLE1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXNOTINTABLE2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXNOTINTABLE3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOOBRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSCALRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSHOLD;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTCFG0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTCFG1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTCFG2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTCFG3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTDONE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTHOLD;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTID00;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTID01;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTID02;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTID03;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTNTRLEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTOVRDEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTPD;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTSTARTED;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTSTROBE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTSTROBEDONE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTSTROBESTARTED;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTTESTOVRDEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSOVRDEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOUTCLK;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOUTCLKFABRIC;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOUTCLKPCS;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOUTCLKSEL0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOUTCLKSEL1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOUTCLKSEL2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPCOMMAALIGNEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPCSRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPD0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPD1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHALIGN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHALIGNDONE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHALIGNEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHDLYPD;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHDLYRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHMONITOR0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHMONITOR1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHMONITOR2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHMONITOR3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHMONITOR4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHOVRDEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHSLIPMONITOR0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHSLIPMONITOR1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHSLIPMONITOR2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHSLIPMONITOR3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHSLIPMONITOR4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPMARESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPMARESETDONE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPOLARITY;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPRBSCNTRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPRBSERR;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPRBSSEL0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPRBSSEL1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPRBSSEL2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXRATE0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXRATE1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXRATE2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXRATEDONE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXRATEMODE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXRESETDONE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSLIDE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSTARTOFSEQ0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSTARTOFSEQ1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSTATUS0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSTATUS1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSTATUS2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSYNCALLIN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSYNCDONE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSYNCIN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSYNCMODE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSYNCOUT;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSYSCLKSEL0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSYSCLKSEL1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXUSERRDY;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXUSRCLK;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXUSRCLK2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXVALID;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_SETERRSTATUS;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_SIGVALIDCLK;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN10;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN11;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN12;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN13;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN14;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN15;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN16;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN17;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN18;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN19;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN5;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN6;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN7;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN8;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN9;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TX8B10BBYPASS0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TX8B10BBYPASS1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TX8B10BBYPASS2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TX8B10BBYPASS3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TX8B10BEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXBUFDIFFCTRL0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXBUFDIFFCTRL1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXBUFDIFFCTRL2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXBUFSTATUS0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXBUFSTATUS1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPMODE0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPMODE1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPMODE2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPMODE3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPVAL0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPVAL1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPVAL2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPVAL3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARISK0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARISK1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARISK2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARISK3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCOMFINISH;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCOMINIT;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCOMSAS;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCOMWAKE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA10;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA11;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA12;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA13;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA14;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA15;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA16;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA17;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA18;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA19;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA20;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA21;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA22;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA23;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA24;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA25;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA26;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA27;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA28;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA29;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA30;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA31;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA5;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA6;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA7;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA8;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA9;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDEEMPH;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDETECTRX;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDIFFCTRL0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDIFFCTRL1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDIFFCTRL2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDIFFCTRL3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDIFFPD;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDLYBYPASS;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDLYEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDLYHOLD;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDLYOVRDEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDLYSRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDLYSRESETDONE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDLYUPDOWN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXELECIDLE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXGEARBOXREADY;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXHEADER0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXHEADER1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXHEADER2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXINHIBIT;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMAINCURSOR0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMAINCURSOR1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMAINCURSOR2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMAINCURSOR3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMAINCURSOR4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMAINCURSOR5;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMAINCURSOR6;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMARGIN0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMARGIN1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMARGIN2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXOUTCLK;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXOUTCLKFABRIC;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXOUTCLKPCS;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXOUTCLKSEL0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXOUTCLKSEL1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXOUTCLKSEL2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPCSRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPD0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPD1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPDELECIDLEMODE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHALIGN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHALIGNDONE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHALIGNEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHDLYPD;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHDLYRESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHDLYTSTCLK;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHINIT;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHINITDONE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHOVRDEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMOVRDEN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMPD;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMSEL;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMSTEPSIZE0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMSTEPSIZE1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMSTEPSIZE2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMSTEPSIZE3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMSTEPSIZE4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPISOPD;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPMARESET;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPMARESETDONE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPOLARITY;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPOSTCURSOR0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPOSTCURSOR1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPOSTCURSOR2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPOSTCURSOR3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPOSTCURSOR4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPOSTCURSORINV;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRBSFORCEERR;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRBSSEL0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRBSSEL1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRBSSEL2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRECURSOR0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRECURSOR1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRECURSOR2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRECURSOR3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRECURSOR4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRECURSORINV;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXRATE0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXRATE1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXRATE2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXRATEDONE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXRATEMODE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXRESETDONE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSEQUENCE0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSEQUENCE1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSEQUENCE2;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSEQUENCE3;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSEQUENCE4;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSEQUENCE5;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSEQUENCE6;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSTARTSEQ;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSWING;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSYNCALLIN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSYNCDONE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSYNCIN;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSYNCMODE;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSYNCOUT;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSYSCLKSEL0;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSYSCLKSEL1;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXUSERRDY;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXUSRCLK;
  wire [0:0] GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXUSRCLK2;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGBYPASSB;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGMONITORENB;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGPDB;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGRCALOVRD0;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGRCALOVRD1;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGRCALOVRD2;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGRCALOVRD3;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGRCALOVRD4;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGRCALOVRDENB;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT0;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT1;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT2;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT3;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT4;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT5;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT6;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT7;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR0;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR1;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR2;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR3;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR4;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR5;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR6;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR7;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPCLK;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI0;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI1;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI10;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI11;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI12;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI13;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI14;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI15;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI2;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI3;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI4;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI5;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI6;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI7;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI8;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI9;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO0;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO1;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO10;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO11;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO12;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO13;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO14;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO15;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO2;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO3;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO4;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO5;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO6;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO7;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO8;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO9;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPEN;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPRDY;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPWE;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_GTREFCLK0;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_GTREFCLK1;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0FBCLKLOST;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0LOCK;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0LOCKDETCLK;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0LOCKEN;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0OUTCLK;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0OUTREFCLK;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0PD;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0REFCLKLOST;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0REFCLKSEL0;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0REFCLKSEL1;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0REFCLKSEL2;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0RESET;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1FBCLKLOST;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1LOCK;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1LOCKDETCLK;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1LOCKEN;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1OUTCLK;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1OUTREFCLK;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1PD;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1REFCLKLOST;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1REFCLKSEL0;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1REFCLKSEL1;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1REFCLKSEL2;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1RESET;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD10;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD11;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD110;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD111;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD112;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD113;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD114;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD115;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD12;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD13;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD14;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD15;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD16;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD17;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD18;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD19;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD20;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD21;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD22;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD23;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD24;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD0;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD1;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD2;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD3;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD4;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD5;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD6;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD7;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT0;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT1;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT10;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT11;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT12;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT13;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT14;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT15;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT2;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT3;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT4;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT5;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT6;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT7;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT8;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT9;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_RCALENB;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_REFCLKOUTMONITOR0;
  wire [0:0] GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_REFCLKOUTMONITOR1;
  wire [0:0] GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y0_CEB;
  wire [0:0] GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y0_O;
  wire [0:0] GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y0_ODIV2;
  wire [0:0] GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y1_CEB;
  wire [0:0] GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y1_O;
  wire [0:0] GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y1_ODIV2;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y11_I;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y3_O;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_O;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_D1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_OQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_T1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_TQ;


  (* KEEP, DONT_TOUCH, BEL = "GTPE2_CHANNEL" *)
  GTPE2_CHANNEL #(
    .ACJTAG_DEBUG_MODE(1'b0),
    .ACJTAG_MODE(1'b0),
    .ACJTAG_RESET(1'b0),
    .ADAPT_CFG0(20'b00000000000000000000),
    .ALIGN_COMMA_DOUBLE("FALSE"),
    .ALIGN_COMMA_ENABLE(10'b0001111111),
    .ALIGN_COMMA_WORD(1),
    .ALIGN_MCOMMA_DET("TRUE"),
    .ALIGN_MCOMMA_VALUE(10'b1010000011),
    .ALIGN_PCOMMA_DET("TRUE"),
    .ALIGN_PCOMMA_VALUE(10'b0101111100),
    .CBCC_DATA_SOURCE_SEL("DECODED"),
    .CFOK_CFG(43'b1001001000000000000000001000000111010000000),
    .CFOK_CFG2(7'b0100000),
    .CFOK_CFG3(7'b0100000),
    .CFOK_CFG4(1'b0),
    .CFOK_CFG5(2'b00),
    .CFOK_CFG6(4'b0000),
    .CHAN_BOND_KEEP_ALIGN("FALSE"),
    .CHAN_BOND_MAX_SKEW(7),
    .CHAN_BOND_SEQ_1_1(10'b0101111100),
    .CHAN_BOND_SEQ_1_2(10'b0000000000),
    .CHAN_BOND_SEQ_1_3(10'b0000000000),
    .CHAN_BOND_SEQ_1_4(10'b0000000000),
    .CHAN_BOND_SEQ_1_ENABLE(4'b1111),
    .CHAN_BOND_SEQ_2_1(10'b0100000000),
    .CHAN_BOND_SEQ_2_2(10'b0100000000),
    .CHAN_BOND_SEQ_2_3(10'b0100000000),
    .CHAN_BOND_SEQ_2_4(10'b0100000000),
    .CHAN_BOND_SEQ_2_ENABLE(4'b1111),
    .CHAN_BOND_SEQ_2_USE("FALSE"),
    .CHAN_BOND_SEQ_LEN(1),
    .CLK_COMMON_SWING(1'b0),
    .CLK_CORRECT_USE("TRUE"),
    .CLK_COR_KEEP_IDLE("FALSE"),
    .CLK_COR_MAX_LAT(20),
    .CLK_COR_MIN_LAT(18),
    .CLK_COR_PRECEDENCE("TRUE"),
    .CLK_COR_REPEAT_WAIT(0),
    .CLK_COR_SEQ_1_1(10'b0100011100),
    .CLK_COR_SEQ_1_2(10'b0000000000),
    .CLK_COR_SEQ_1_3(10'b0000000000),
    .CLK_COR_SEQ_1_4(10'b0000000000),
    .CLK_COR_SEQ_1_ENABLE(4'b1111),
    .CLK_COR_SEQ_2_1(10'b0100000000),
    .CLK_COR_SEQ_2_2(10'b0100000000),
    .CLK_COR_SEQ_2_3(10'b0100000000),
    .CLK_COR_SEQ_2_4(10'b0100000000),
    .CLK_COR_SEQ_2_ENABLE(4'b1111),
    .CLK_COR_SEQ_2_USE("FALSE"),
    .CLK_COR_SEQ_LEN(1),
    .DEC_MCOMMA_DETECT("TRUE"),
    .DEC_PCOMMA_DETECT("TRUE"),
    .DEC_VALID_COMMA_ONLY("TRUE"),
    .DMONITOR_CFG(24'b000000000000101000000000),
    .ES_CLK_PHASE_SEL(1'b0),
    .ES_CONTROL(6'b000000),
    .ES_ERRDET_EN("FALSE"),
    .ES_EYE_SCAN_EN("FALSE"),
    .ES_HORZ_OFFSET(12'b000000010000),
    .ES_PMA_CFG(10'b0000000000),
    .ES_PRESCALE(5'b00000),
    .ES_QUALIFIER(80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000),
    .ES_QUAL_MASK(80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000),
    .ES_SDATA_MASK(80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000),
    .ES_VERT_OFFSET(9'b000000000),
    .FTS_DESKEW_SEQ_ENABLE(4'b1111),
    .FTS_LANE_DESKEW_CFG(4'b1111),
    .FTS_LANE_DESKEW_EN("FALSE"),
    .GEARBOX_MODE(3'b000),
    .IS_CLKRSVD0_INVERTED(1),
    .IS_CLKRSVD1_INVERTED(1),
    .IS_DMONITORCLK_INVERTED(1),
    .IS_RXUSRCLK2_INVERTED(1),
    .IS_RXUSRCLK_INVERTED(1),
    .IS_SIGVALIDCLK_INVERTED(1),
    .IS_TXPHDLYTSTCLK_INVERTED(1),
    .IS_TXUSRCLK2_INVERTED(1),
    .IS_TXUSRCLK_INVERTED(1),
    .LOOPBACK_CFG(1'b0),
    .OUTREFCLK_SEL_INV(2'b11),
    .PCS_PCIE_EN("FALSE"),
    .PCS_RSVD_ATTR(48'b000000000000000000000000000000000000000000000000),
    .PD_TRANS_TIME_FROM_P2(12'b000000111100),
    .PD_TRANS_TIME_NONE_P2(8'b00011001),
    .PD_TRANS_TIME_TO_P2(8'b01100100),
    .PMA_LOOPBACK_CFG(1'b0),
    .PMA_RSV(32'b00000000000000000000001100110011),
    .PMA_RSV2(32'b00000000000000000010000001010000),
    .PMA_RSV3(2'b00),
    .PMA_RSV4(4'b0000),
    .PMA_RSV5(1'b0),
    .PMA_RSV6(1'b0),
    .PMA_RSV7(1'b0),
    .RXBUFRESET_TIME(5'b00001),
    .RXBUF_ADDR_MODE("FULL"),
    .RXBUF_EIDLE_HI_CNT(4'b1000),
    .RXBUF_EIDLE_LO_CNT(4'b0000),
    .RXBUF_EN("TRUE"),
    .RXBUF_RESET_ON_CB_CHANGE("TRUE"),
    .RXBUF_RESET_ON_COMMAALIGN("FALSE"),
    .RXBUF_RESET_ON_EIDLE("FALSE"),
    .RXBUF_RESET_ON_RATE_CHANGE("TRUE"),
    .RXBUF_THRESH_OVFLW(61),
    .RXBUF_THRESH_OVRD("FALSE"),
    .RXBUF_THRESH_UNDFLW(4),
    .RXCDRFREQRESET_TIME(5'b00001),
    .RXCDRPHRESET_TIME(5'b00001),
    .RXCDR_CFG(83'b00000000000000000010000011111111110010000000110000000000001000001000001000000010000),
    .RXCDR_FR_RESET_ON_EIDLE(1'b0),
    .RXCDR_HOLD_DURING_EIDLE(1'b0),
    .RXCDR_LOCK_CFG(6'b001001),
    .RXCDR_PH_RESET_ON_EIDLE(1'b0),
    .RXDLY_CFG(16'b0000000000010000),
    .RXDLY_LCFG(9'b000100000),
    .RXDLY_TAP_CFG(16'b0000000000000000),
    .RXGEARBOX_EN("FALSE"),
    .RXISCANRESET_TIME(5'b00001),
    .RXLPMRESET_TIME(7'b0001111),
    .RXLPM_BIAS_STARTUP_DISABLE(1'b0),
    .RXLPM_CFG(4'b0110),
    .RXLPM_CFG1(1'b0),
    .RXLPM_CM_CFG(1'b0),
    .RXLPM_GC_CFG(9'b111100010),
    .RXLPM_GC_CFG2(3'b001),
    .RXLPM_HF_CFG(14'b00001111110000),
    .RXLPM_HF_CFG2(5'b01010),
    .RXLPM_HF_CFG3(4'b0000),
    .RXLPM_HOLD_DURING_EIDLE(1'b0),
    .RXLPM_INCM_CFG(1'b0),
    .RXLPM_IPCM_CFG(1'b0),
    .RXLPM_LF_CFG(18'b000000001111110000),
    .RXLPM_LF_CFG2(5'b01010),
    .RXLPM_OSINT_CFG(3'b100),
    .RXOOB_CFG(7'b0000110),
    .RXOOB_CLK_CFG("PMA"),
    .RXOSCALRESET_TIME(5'b00011),
    .RXOSCALRESET_TIMEOUT(5'b00000),
    .RXOUT_DIV(2),
    .RXPCSRESET_TIME(5'b00001),
    .RXPHDLY_CFG(24'b000010000100000000000000),
    .RXPH_CFG(24'b110000000000000000000010),
    .RXPH_MONITOR_SEL(5'b00000),
    .RXPI_CFG0(3'b000),
    .RXPI_CFG1(1'b0),
    .RXPI_CFG2(1'b0),
    .RXPMARESET_TIME(5'b00011),
    .RXPRBS_ERR_LOOPBACK(1'b0),
    .RXSLIDE_AUTO_WAIT(7),
    .RXSLIDE_MODE("OFF"),
    .RXSYNC_MULTILANE(1'b0),
    .RXSYNC_OVRD(1'b0),
    .RXSYNC_SKIP_DA(1'b0),
    .RX_BIAS_CFG(16'b0000111100110011),
    .RX_BUFFER_CFG(6'b000000),
    .RX_CLK25_DIV(7),
    .RX_CLKMUX_EN(1'b1),
    .RX_CM_SEL(2'b11),
    .RX_CM_TRIM(4'b0100),
    .RX_DATA_WIDTH(20),
    .RX_DDI_SEL(6'b000000),
    .RX_DEBUG_CFG(14'b00000000000000),
    .RX_DEFER_RESET_BUF_EN("TRUE"),
    .RX_DISPERR_SEQ_MATCH("TRUE"),
    .RX_OS_CFG(13'b0001111110000),
    .RX_SIG_VALID_DLY(10),
    .RX_XCLK_SEL("RXREC"),
    .SAS_MAX_COM(64),
    .SAS_MIN_COM(36),
    .SATA_BURST_SEQ_LEN(4'b1111),
    .SATA_BURST_VAL(3'b100),
    .SATA_EIDLE_VAL(3'b100),
    .SATA_MAX_BURST(8),
    .SATA_MAX_INIT(21),
    .SATA_MAX_WAKE(7),
    .SATA_MIN_BURST(4),
    .SATA_MIN_INIT(12),
    .SATA_MIN_WAKE(4),
    .SATA_PLL_CFG("VCO_3000MHZ"),
    .SHOW_REALIGN_COMMA("TRUE"),
    .TERM_RCAL_CFG(15'b100001000010000),
    .TERM_RCAL_OVRD(3'b000),
    .TRANS_TIME_RATE(8'b00001110),
    .TST_RSV(32'b00000000000000000000000000000000),
    .TXBUF_EN("TRUE"),
    .TXBUF_RESET_ON_RATE_CHANGE("FALSE"),
    .TXDLY_CFG(16'b0000000000010000),
    .TXDLY_LCFG(9'b000100000),
    .TXDLY_TAP_CFG(16'b0000000000000000),
    .TXGEARBOX_EN("FALSE"),
    .TXOOB_CFG(1'b0),
    .TXOUT_DIV(2),
    .TXPCSRESET_TIME(5'b00001),
    .TXPHDLY_CFG(24'b000010000100000000000000),
    .TXPH_CFG(16'b0000010000000000),
    .TXPH_MONITOR_SEL(5'b00000),
    .TXPI_CFG0(2'b00),
    .TXPI_CFG1(2'b00),
    .TXPI_CFG2(2'b00),
    .TXPI_CFG3(1'b0),
    .TXPI_CFG4(1'b0),
    .TXPI_CFG5(3'b000),
    .TXPI_GREY_SEL(1'b0),
    .TXPI_INVSTROBE_SEL(1'b0),
    .TXPI_PPMCLK_SEL("TXUSRCLK2"),
    .TXPI_PPM_CFG(8'b00000000),
    .TXPI_SYNFREQ_PPM(3'b000),
    .TXPMARESET_TIME(5'b00001),
    .TXSYNC_MULTILANE(1'b0),
    .TXSYNC_OVRD(1'b0),
    .TXSYNC_SKIP_DA(1'b0),
    .TX_CLK25_DIV(7),
    .TX_CLKMUX_EN(1'b1),
    .TX_DATA_WIDTH(20),
    .TX_DEEMPH0(6'b000000),
    .TX_DEEMPH1(6'b000000),
    .TX_DRIVE_MODE("DIRECT"),
    .TX_EIDLE_ASSERT_DELAY(3'b110),
    .TX_EIDLE_DEASSERT_DELAY(3'b100),
    .TX_LOOPBACK_DRIVE_HIZ("FALSE"),
    .TX_MAINCURSOR_SEL(1'b0),
    .TX_MARGIN_FULL_0(7'b1001110),
    .TX_MARGIN_FULL_1(7'b1001001),
    .TX_MARGIN_FULL_2(7'b1000101),
    .TX_MARGIN_FULL_3(7'b1000010),
    .TX_MARGIN_FULL_4(7'b1000000),
    .TX_MARGIN_LOW_0(7'b1000110),
    .TX_MARGIN_LOW_1(7'b1000100),
    .TX_MARGIN_LOW_2(7'b1000010),
    .TX_MARGIN_LOW_3(7'b1000000),
    .TX_MARGIN_LOW_4(7'b1000000),
    .TX_PREDRIVER_MODE(1'b0),
    .TX_RXDETECT_CFG(14'b01100000110010),
    .TX_RXDETECT_REF(3'b100),
    .TX_XCLK_SEL("TXUSR"),
    .UCODEER_CLR(1'b0),
    .USE_PCS_CLK_PHASE_SEL(1'b0)
  ) GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTPE2_CHANNEL (
.CFGRESET(1'b0),
.CLKRSVD0(1'b1),
.CLKRSVD1(1'b1),
.DMONFIFORESET(1'b0),
.DMONITORCLK(1'b1),
.DMONITOROUT({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT14, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT13, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT12, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT11, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT10, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT9, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT8, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT7, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT6, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT5, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT4, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT3, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT2, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITOROUT0}),
.DRPADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b1}),
.DRPCLK(1'b1),
.DRPDI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1}),
.DRPDO({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO15, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO14, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO13, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO12, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO11, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO10, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO9, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO8, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO7, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO6, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO5, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO4, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO3, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO2, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDO0}),
.DRPEN(LIOB33_X0Y11_IOB_X0Y11_I),
.DRPRDY(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPRDY),
.DRPWE(LIOB33_X0Y11_IOB_X0Y11_I),
.EYESCANDATAERROR(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_EYESCANDATAERROR),
.EYESCANMODE(1'b0),
.EYESCANRESET(1'b0),
.EYESCANTRIGGER(1'b0),
.GTPRXN(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_IPAD_RX_N),
.GTPRXP(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_IPAD_RX_P),
.GTPTXN(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_OPAD_TX_N),
.GTPTXP(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_OPAD_TX_P),
.GTRESETSEL(1'b0),
.GTRSVD({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.GTRXRESET(1'b0),
.GTTXRESET(1'b0),
.LOOPBACK({1'b0, 1'b0, 1'b0}),
.PCSRSVDIN({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.PCSRSVDOUT({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT15, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT14, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT13, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT12, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT11, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT10, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT9, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT8, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT7, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT6, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT5, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT4, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT3, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT2, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDOUT0}),
.PHYSTATUS(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PHYSTATUS),
.PMARSVDIN0(1'b0),
.PMARSVDIN1(1'b0),
.PMARSVDIN2(1'b0),
.PMARSVDIN3(1'b0),
.PMARSVDIN4(1'b0),
.PMARSVDOUT0(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PMARSVDOUT0),
.PMARSVDOUT1(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PMARSVDOUT1),
.RESETOVRD(1'b0),
.RX8B10BEN(1'b0),
.RXADAPTSELTEST({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.RXBUFRESET(1'b0),
.RXBUFSTATUS({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXBUFSTATUS2, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXBUFSTATUS1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXBUFSTATUS0}),
.RXBYTEISALIGNED(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXBYTEISALIGNED),
.RXBYTEREALIGN(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXBYTEREALIGN),
.RXCDRFREQRESET(1'b0),
.RXCDRHOLD(1'b0),
.RXCDRLOCK(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCDRLOCK),
.RXCDROVRDEN(1'b0),
.RXCDRRESET(1'b0),
.RXCDRRESETRSV(1'b0),
.RXCHANBONDSEQ(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHANBONDSEQ),
.RXCHANISALIGNED(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHANISALIGNED),
.RXCHANREALIGN(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHANREALIGN),
.RXCHARISCOMMA({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISCOMMA3, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISCOMMA2, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISCOMMA1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISCOMMA0}),
.RXCHARISK({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISK3, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISK2, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISK1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHARISK0}),
.RXCHBONDEN(1'b0),
.RXCHBONDI({1'b0, 1'b0, 1'b0, 1'b0}),
.RXCHBONDLEVEL({1'b0, 1'b0, 1'b0}),
.RXCHBONDMASTER(1'b0),
.RXCHBONDO({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDO3, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDO2, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDO1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDO0}),
.RXCHBONDSLAVE(1'b0),
.RXCLKCORCNT({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCLKCORCNT1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCLKCORCNT0}),
.RXCOMINITDET(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCOMINITDET),
.RXCOMMADET(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCOMMADET),
.RXCOMMADETEN(1'b0),
.RXCOMSASDET(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCOMSASDET),
.RXCOMWAKEDET(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCOMWAKEDET),
.RXDATA({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA31, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA30, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA29, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA28, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA27, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA26, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA25, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA24, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA23, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA22, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA21, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA20, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA19, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA18, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA17, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA16, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA15, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA14, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA13, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA12, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA11, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA10, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA9, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA8, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA7, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA6, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA5, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA4, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA3, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA2, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATA0}),
.RXDATAVALID({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATAVALID1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDATAVALID0}),
.RXDDIEN(1'b0),
.RXDFEXYDEN(1'b0),
.RXDISPERR({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDISPERR3, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDISPERR2, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDISPERR1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDISPERR0}),
.RXDLYBYPASS(1'b0),
.RXDLYEN(1'b0),
.RXDLYOVRDEN(1'b0),
.RXDLYSRESET(1'b0),
.RXDLYSRESETDONE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDLYSRESETDONE),
.RXELECIDLE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXELECIDLE),
.RXELECIDLEMODE({1'b0, 1'b0}),
.RXGEARBOXSLIP(1'b0),
.RXHEADER({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXHEADER2, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXHEADER1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXHEADER0}),
.RXHEADERVALID(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXHEADERVALID),
.RXLPMHFHOLD(1'b0),
.RXLPMHFOVRDEN(1'b0),
.RXLPMLFHOLD(1'b0),
.RXLPMLFOVRDEN(1'b0),
.RXLPMOSINTNTRLEN(1'b0),
.RXLPMRESET(1'b0),
.RXMCOMMAALIGNEN(1'b0),
.RXNOTINTABLE({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXNOTINTABLE3, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXNOTINTABLE2, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXNOTINTABLE1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXNOTINTABLE0}),
.RXOOBRESET(1'b0),
.RXOSCALRESET(1'b0),
.RXOSHOLD(1'b0),
.RXOSINTCFG({1'b0, 1'b0, 1'b0, 1'b0}),
.RXOSINTDONE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTDONE),
.RXOSINTEN(1'b0),
.RXOSINTHOLD(1'b0),
.RXOSINTID0({1'b0, 1'b0, 1'b0, 1'b0}),
.RXOSINTNTRLEN(1'b0),
.RXOSINTOVRDEN(1'b0),
.RXOSINTPD(1'b0),
.RXOSINTSTARTED(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTSTARTED),
.RXOSINTSTROBE(1'b0),
.RXOSINTSTROBEDONE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTSTROBEDONE),
.RXOSINTSTROBESTARTED(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTSTROBESTARTED),
.RXOSINTTESTOVRDEN(1'b0),
.RXOSOVRDEN(1'b0),
.RXOUTCLK(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOUTCLK),
.RXOUTCLKFABRIC(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOUTCLKFABRIC),
.RXOUTCLKPCS(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOUTCLKPCS),
.RXOUTCLKSEL({1'b0, 1'b0, 1'b0}),
.RXPCOMMAALIGNEN(1'b0),
.RXPCSRESET(1'b0),
.RXPD({1'b0, 1'b0}),
.RXPHALIGN(1'b0),
.RXPHALIGNDONE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHALIGNDONE),
.RXPHALIGNEN(1'b0),
.RXPHDLYPD(1'b0),
.RXPHDLYRESET(1'b0),
.RXPHMONITOR({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHMONITOR4, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHMONITOR3, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHMONITOR2, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHMONITOR1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHMONITOR0}),
.RXPHOVRDEN(1'b0),
.RXPHSLIPMONITOR({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHSLIPMONITOR4, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHSLIPMONITOR3, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHSLIPMONITOR2, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHSLIPMONITOR1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHSLIPMONITOR0}),
.RXPMARESET(1'b0),
.RXPMARESETDONE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPMARESETDONE),
.RXPOLARITY(1'b0),
.RXPRBSCNTRESET(1'b0),
.RXPRBSERR(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPRBSERR),
.RXPRBSSEL({1'b0, 1'b0, 1'b0}),
.RXRATE({1'b0, 1'b0, 1'b0}),
.RXRATEDONE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXRATEDONE),
.RXRATEMODE(1'b0),
.RXRESETDONE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXRESETDONE),
.RXSLIDE(1'b0),
.RXSTARTOFSEQ({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSTARTOFSEQ1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSTARTOFSEQ0}),
.RXSTATUS({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSTATUS2, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSTATUS1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSTATUS0}),
.RXSYNCALLIN(1'b0),
.RXSYNCDONE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSYNCDONE),
.RXSYNCIN(1'b0),
.RXSYNCMODE(1'b0),
.RXSYNCOUT(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSYNCOUT),
.RXSYSCLKSEL({1'b0, 1'b0}),
.RXUSERRDY(1'b0),
.RXUSRCLK(1'b1),
.RXUSRCLK2(1'b1),
.RXVALID(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXVALID),
.SETERRSTATUS(1'b0),
.SIGVALIDCLK(1'b1),
.TSTIN({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.TX8B10BBYPASS({1'b0, 1'b0, 1'b0, 1'b0}),
.TX8B10BEN(1'b0),
.TXBUFDIFFCTRL({1'b0, 1'b0, 1'b0}),
.TXBUFSTATUS({GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXBUFSTATUS1, GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXBUFSTATUS0}),
.TXCHARDISPMODE({1'b0, 1'b0, 1'b0, 1'b0}),
.TXCHARDISPVAL({1'b0, 1'b0, 1'b0, 1'b0}),
.TXCHARISK({1'b0, 1'b0, 1'b0, 1'b0}),
.TXCOMFINISH(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCOMFINISH),
.TXCOMINIT(1'b0),
.TXCOMSAS(1'b0),
.TXCOMWAKE(1'b0),
.TXDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.TXDEEMPH(1'b0),
.TXDETECTRX(1'b0),
.TXDIFFCTRL({1'b0, 1'b0, 1'b0, 1'b0}),
.TXDIFFPD(1'b0),
.TXDLYBYPASS(1'b0),
.TXDLYEN(1'b0),
.TXDLYHOLD(1'b0),
.TXDLYOVRDEN(1'b0),
.TXDLYSRESET(1'b0),
.TXDLYSRESETDONE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDLYSRESETDONE),
.TXDLYUPDOWN(1'b0),
.TXELECIDLE(1'b0),
.TXGEARBOXREADY(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXGEARBOXREADY),
.TXHEADER({1'b0, 1'b0, 1'b0}),
.TXINHIBIT(1'b0),
.TXMAINCURSOR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.TXMARGIN({1'b0, 1'b0, 1'b0}),
.TXOUTCLK(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXOUTCLK),
.TXOUTCLKFABRIC(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXOUTCLKFABRIC),
.TXOUTCLKPCS(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXOUTCLKPCS),
.TXOUTCLKSEL({1'b0, 1'b0, 1'b0}),
.TXPCSRESET(1'b0),
.TXPD({1'b0, 1'b0}),
.TXPDELECIDLEMODE(1'b0),
.TXPHALIGN(1'b0),
.TXPHALIGNDONE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHALIGNDONE),
.TXPHALIGNEN(1'b0),
.TXPHDLYPD(1'b0),
.TXPHDLYRESET(1'b0),
.TXPHDLYTSTCLK(1'b1),
.TXPHINIT(1'b0),
.TXPHINITDONE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHINITDONE),
.TXPHOVRDEN(1'b0),
.TXPIPPMEN(1'b0),
.TXPIPPMOVRDEN(1'b0),
.TXPIPPMPD(1'b0),
.TXPIPPMSEL(1'b0),
.TXPIPPMSTEPSIZE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.TXPISOPD(1'b0),
.TXPMARESET(1'b0),
.TXPMARESETDONE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPMARESETDONE),
.TXPOLARITY(1'b0),
.TXPOSTCURSOR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.TXPOSTCURSORINV(1'b0),
.TXPRBSFORCEERR(1'b0),
.TXPRBSSEL({1'b0, 1'b0, 1'b0}),
.TXPRECURSOR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.TXPRECURSORINV(1'b0),
.TXRATE({1'b0, 1'b0, 1'b0}),
.TXRATEDONE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXRATEDONE),
.TXRATEMODE(1'b0),
.TXRESETDONE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXRESETDONE),
.TXSEQUENCE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.TXSTARTSEQ(1'b0),
.TXSWING(1'b0),
.TXSYNCALLIN(1'b0),
.TXSYNCDONE(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSYNCDONE),
.TXSYNCIN(1'b0),
.TXSYNCMODE(1'b0),
.TXSYNCOUT(GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSYNCOUT),
.TXSYSCLKSEL({1'b0, 1'b0}),
.TXUSERRDY(1'b0),
.TXUSRCLK(1'b1),
.TXUSRCLK2(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "IBUFDS_GTE2" *)
  IBUFDS_GTE2 #(
    .CLKCM_CFG("TRUE"),
    .CLKRCV_TRST("TRUE")
  ) GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y0_IBUFDS_GTE2 (
.CEB(1'b0),
.I(GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y0_IPAD_P),
.IB(GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y0_IPAD_N),
.O(GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y0_O),
.ODIV2(GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y0_ODIV2)
  );


  (* KEEP, DONT_TOUCH, BEL = "IBUFDS_GTE2" *)
  IBUFDS_GTE2 #(
    .CLKCM_CFG("TRUE"),
    .CLKRCV_TRST("TRUE")
  ) GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y1_IBUFDS_GTE2 (
.CEB(1'b0),
.I(GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y1_IPAD_P),
.IB(GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y1_IPAD_N),
.O(GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y1_O),
.ODIV2(GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y1_ODIV2)
  );


  (* KEEP, DONT_TOUCH, BEL = "GTPE2_COMMON" *)
  GTPE2_COMMON #(
    .BIAS_CFG(64'b0000000000000000000000000000000000000000000000000000000000000000),
    .COMMON_CFG(32'b00000000000000000000000000000000),
    .IS_DRPCLK_INVERTED(1),
    .IS_PLL0LOCKDETCLK_INVERTED(1),
    .IS_PLL1LOCKDETCLK_INVERTED(1),
    .PLL0_CFG(27'b000000111110000001111011100),
    .PLL0_DMON_CFG(1'b0),
    .PLL0_FBDIV(5),
    .PLL0_FBDIV_45(4),
    .PLL0_INIT_CFG(24'b000000000000000000011110),
    .PLL0_LOCK_CFG(9'b111101000),
    .PLL0_REFCLK_DIV(1),
    .PLL1_CFG(27'b000000111110000001111011100),
    .PLL1_DMON_CFG(1'b0),
    .PLL1_FBDIV(4),
    .PLL1_FBDIV_45(5),
    .PLL1_INIT_CFG(24'b000000000000000000011110),
    .PLL1_LOCK_CFG(9'b111101000),
    .PLL1_REFCLK_DIV(1),
    .PLL_CLKOUT_CFG(8'b00000000),
    .RSVD_ATTR0(16'b0000000000000000),
    .RSVD_ATTR1(16'b0000000000000000)
  ) GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_GTPE2_COMMON (
.BGBYPASSB(1'b1),
.BGMONITORENB(LIOB33_X0Y11_IOB_X0Y11_I),
.BGPDB(1'b1),
.BGRCALOVRD({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.BGRCALOVRDENB(1'b0),
.DMONITOROUT({GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT7, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT6, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT5, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT4, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT3, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT2, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT1, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DMONITOROUT0}),
.DRPADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.DRPCLK(1'b1),
.DRPDI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.DRPDO({GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO15, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO14, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO13, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO12, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO11, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO10, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO9, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO8, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO7, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO6, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO5, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO4, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO3, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO2, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO1, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDO0}),
.DRPEN(1'b0),
.DRPRDY(GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPRDY),
.DRPWE(1'b0),
.GTREFCLK0(GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y0_O),
.GTREFCLK1(GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y1_O),
.PLL0FBCLKLOST(GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0FBCLKLOST),
.PLL0LOCK(GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0LOCK),
.PLL0LOCKDETCLK(1'b1),
.PLL0LOCKEN(1'b1),
.PLL0OUTCLK(GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0OUTCLK),
.PLL0OUTREFCLK(GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0OUTREFCLK),
.PLL0PD(1'b0),
.PLL0REFCLKLOST(GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0REFCLKLOST),
.PLL0REFCLKSEL({1'b0, 1'b0, 1'b1}),
.PLL0RESET(1'b0),
.PLL1FBCLKLOST(GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1FBCLKLOST),
.PLL1LOCK(GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1LOCK),
.PLL1LOCKDETCLK(1'b1),
.PLL1LOCKEN(1'b0),
.PLL1OUTCLK(GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1OUTCLK),
.PLL1OUTREFCLK(GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1OUTREFCLK),
.PLL1PD(1'b1),
.PLL1REFCLKLOST(GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1REFCLKLOST),
.PLL1REFCLKSEL({1'b0, 1'b0, 1'b0}),
.PLL1RESET(1'b0),
.PLLRSVD1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.PLLRSVD2({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}),
.PMARSVD({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.PMARSVDOUT({GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT15, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT14, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT13, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT12, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT11, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT10, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT9, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT8, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT7, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT6, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT5, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT4, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT3, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT2, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT1, GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVDOUT0}),
.RCALENB(1'b1),
.REFCLKOUTMONITOR0(GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_REFCLKOUTMONITOR0),
.REFCLKOUTMONITOR1(GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_REFCLKOUTMONITOR1)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y3_IOB_X0Y3_OBUF (
.I(GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_REFCLKOUTMONITOR0),
.O(test_out)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y11_IOB_X0Y11_IBUF (
.I(test_in),
.O(LIOB33_X0Y11_IOB_X0Y11_I)
  );
  assign LIOI3_X0Y3_OLOGIC_X0Y3_OQ = GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_REFCLKOUTMONITOR0;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_TQ = 1'b1;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_O = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOB33_X0Y3_IOB_X0Y3_O = GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_REFCLKOUTMONITOR0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD0 = 1'b0;
  assign GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y0_CEB = 1'b0;
  assign GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y1_CEB = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR7 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPCLK = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI0 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI7 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI8 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI9 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI10 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI11 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD4 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI12 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_CFGRESET = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_CLKRSVD0 = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_CLKRSVD1 = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONFIFORESET = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DMONITORCLK = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI13 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI15 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR0 = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR4 = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR5 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR6 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR7 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPADDR8 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPCLK = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI0 = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI4 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI5 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI6 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI7 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI8 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI9 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI10 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI11 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI12 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI13 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI14 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPDI15 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPEN = LIOB33_X0Y11_IOB_X0Y11_I;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_DRPWE = LIOB33_X0Y11_IOB_X0Y11_I;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_EYESCANMODE = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_EYESCANRESET = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_EYESCANTRIGGER = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRESETSEL = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD4 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD5 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD6 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD7 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD8 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD9 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD10 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD11 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD12 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD13 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD14 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRSVD15 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTRXRESET = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_GTTXRESET = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_LOOPBACK0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_LOOPBACK1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_LOOPBACK2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN4 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN5 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN6 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN7 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN8 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN9 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN10 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN11 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN12 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN13 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN14 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PCSRSVDIN15 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PMARSVDIN0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PMARSVDIN1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PMARSVDIN2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PMARSVDIN3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_PMARSVDIN4 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RESETOVRD = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RX8B10BEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST4 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST5 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST6 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST7 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST8 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST9 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST10 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST11 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST12 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXADAPTSELTEST13 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXBUFRESET = 1'b0;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_D1 = GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_REFCLKOUTMONITOR0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCDRFREQRESET = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCDRHOLD = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCDROVRDEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCDRRESET = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCDRRESETRSV = 1'b0;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_T1 = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDI0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDI1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDI2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDI3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDLEVEL0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDLEVEL1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDLEVEL2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDMASTER = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCHBONDSLAVE = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXCOMMADETEN = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGBYPASSB = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGMONITORENB = LIOB33_X0Y11_IOB_X0Y11_I;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGPDB = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGRCALOVRD0 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGRCALOVRD1 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGRCALOVRD2 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGRCALOVRD3 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGRCALOVRD4 = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDDIEN = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_BGRCALOVRDENB = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDFEXYDEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDLYBYPASS = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDLYEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDLYOVRDEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXDLYSRESET = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR0 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR1 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXELECIDLEMODE0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXELECIDLEMODE1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXGEARBOXSLIP = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR3 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR4 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR5 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPADDR6 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXLPMHFHOLD = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXLPMHFOVRDEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXLPMLFHOLD = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXLPMLFOVRDEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXLPMOSINTNTRLEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXLPMRESET = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXMCOMMAALIGNEN = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI1 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI2 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI3 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI4 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI5 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI6 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOOBRESET = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSCALRESET = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSHOLD = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTCFG0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTCFG1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTCFG2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTCFG3 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPDI14 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTHOLD = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTID00 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTID01 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTID02 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTID03 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTNTRLEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTOVRDEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTPD = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTSTROBE = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_DRPWE = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSINTTESTOVRDEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOSOVRDEN = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_GTREFCLK0 = GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y0_O;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_GTREFCLK1 = GTP_COMMON_X97Y127_IBUFDS_GTE2_X0Y1_O;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOUTCLKSEL0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOUTCLKSEL1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXOUTCLKSEL2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPCOMMAALIGNEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPCSRESET = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPD0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPD1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHALIGN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHALIGNEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHDLYPD = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHDLYRESET = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0LOCKDETCLK = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0LOCKEN = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0PD = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0REFCLKSEL0 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0REFCLKSEL1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPHOVRDEN = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0REFCLKSEL2 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL0RESET = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1LOCKDETCLK = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1LOCKEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPMARESET = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1PD = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPOLARITY = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPRBSCNTRESET = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1REFCLKSEL0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPRBSSEL0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPRBSSEL1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXPRBSSEL2 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1REFCLKSEL1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXRATE0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXRATE1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXRATE2 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1REFCLKSEL2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXRATEMODE = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLL1RESET = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSLIDE = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD10 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD11 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD12 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD13 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD14 = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSYNCALLIN = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD15 = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSYNCIN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSYNCMODE = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD16 = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSYSCLKSEL0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXSYSCLKSEL1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXUSERRDY = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXUSRCLK = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_RXUSRCLK2 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD19 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD20 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD21 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD22 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD23 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD24 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD110 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD111 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD112 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD113 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD114 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD115 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD17 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD1 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD2 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_SETERRSTATUS = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_SIGVALIDCLK = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PLLRSVD18 = 1'b1;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD7 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN4 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN5 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN6 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN7 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN8 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN9 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN10 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN11 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN12 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN13 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN14 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN15 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN16 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN17 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN18 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TSTIN19 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_RCALENB = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TX8B10BBYPASS0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TX8B10BBYPASS1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TX8B10BBYPASS2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TX8B10BBYPASS3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TX8B10BEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXBUFDIFFCTRL0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXBUFDIFFCTRL1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXBUFDIFFCTRL2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPMODE0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPMODE1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPMODE2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPMODE3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPVAL0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPVAL1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPVAL2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARDISPVAL3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARISK0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARISK1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARISK2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCHARISK3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCOMINIT = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCOMSAS = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXCOMWAKE = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA4 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA5 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA6 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA7 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA8 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA9 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA10 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA11 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA12 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA13 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA14 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA15 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA16 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA17 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA18 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA19 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA20 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA21 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA22 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA23 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA24 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA25 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA26 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA27 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA28 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA29 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA30 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDATA31 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDEEMPH = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDETECTRX = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDIFFCTRL0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDIFFCTRL1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDIFFCTRL2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDIFFCTRL3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDIFFPD = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDLYBYPASS = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDLYEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDLYHOLD = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDLYOVRDEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDLYSRESET = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD5 = 1'b0;
  assign GTP_COMMON_X97Y127_GTPE2_COMMON_X0Y0_PMARSVD6 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXDLYUPDOWN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXELECIDLE = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXHEADER0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXHEADER1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXHEADER2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXINHIBIT = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMAINCURSOR0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMAINCURSOR1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMAINCURSOR2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMAINCURSOR3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMAINCURSOR4 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMAINCURSOR5 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMAINCURSOR6 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMARGIN0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMARGIN1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXMARGIN2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXOUTCLKSEL0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXOUTCLKSEL1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXOUTCLKSEL2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPCSRESET = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPD0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPD1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPDELECIDLEMODE = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHALIGN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHALIGNEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHDLYPD = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHDLYRESET = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHDLYTSTCLK = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHINIT = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPHOVRDEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMOVRDEN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMPD = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMSEL = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMSTEPSIZE0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMSTEPSIZE1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMSTEPSIZE2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMSTEPSIZE3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPIPPMSTEPSIZE4 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPISOPD = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPMARESET = 1'b0;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_D = LIOB33_X0Y11_IOB_X0Y11_I;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPOLARITY = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPOSTCURSOR0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPOSTCURSOR1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPOSTCURSOR2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPOSTCURSOR3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPOSTCURSOR4 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPOSTCURSORINV = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRBSFORCEERR = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRBSSEL0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRBSSEL1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRBSSEL2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRECURSOR0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRECURSOR1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRECURSOR2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRECURSOR3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRECURSOR4 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXPRECURSORINV = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXRATE0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXRATE1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXRATE2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXRATEMODE = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSEQUENCE0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSEQUENCE1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSEQUENCE2 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSEQUENCE3 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSEQUENCE4 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSEQUENCE5 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSEQUENCE6 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSTARTSEQ = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSWING = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSYNCALLIN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSYNCIN = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSYNCMODE = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSYSCLKSEL0 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXSYSCLKSEL1 = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXUSERRDY = 1'b0;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXUSRCLK = 1'b1;
  assign GTP_CHANNEL_0_X97Y110_GTPE2_CHANNEL_X0Y0_TXUSRCLK2 = 1'b1;
endmodule
