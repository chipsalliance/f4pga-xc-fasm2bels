module top(
  input i_ce,
  input i_clk,
  input i_clkb,
  input i_rst,
  input [35:0] io,
  output o_q1,
  output o_q2
  );
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_A;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_A1;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_A2;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_A3;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_A4;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_A5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_A6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_AMUX;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_AO5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_AO6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_A_CY;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_A_XOR;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_B;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_B1;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_B2;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_B3;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_B4;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_B5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_B6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_BMUX;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_BO5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_BO6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_B_CY;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_B_XOR;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_C;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_C1;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_C2;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_C3;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_C4;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_C5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_C6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_CMUX;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_CO5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_CO6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_C_CY;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_C_XOR;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_D;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_D1;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_D2;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_D3;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_D4;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_D5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_D6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_DMUX;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_DO5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_DO6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_D_CY;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X0Y22_D_XOR;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_A;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_A1;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_A2;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_A3;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_A4;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_A5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_A6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_AO5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_AO6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_A_CY;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_A_XOR;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_B;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_B1;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_B2;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_B3;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_B4;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_B5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_B6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_BO5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_BO6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_B_CY;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_B_XOR;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_C;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_C1;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_C2;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_C3;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_C4;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_C5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_C6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_CO5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_CO6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_C_CY;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_C_XOR;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_D;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_D1;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_D2;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_D3;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_D4;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_D5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_D6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_DO5;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_DO6;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_D_CY;
  wire [0:0] CLBLL_L_X2Y22_SLICE_X1Y22_D_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_AMUX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_AO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_AO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_BMUX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_BO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_BO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_CMUX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_CO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_CO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_DMUX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_DO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_DO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_AMUX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_AO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_AO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_BMUX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_BO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_BO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_CMUX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_CO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_CO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_DMUX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_DO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_DO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_AMUX;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_AO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_AO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_BMUX;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_BO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_BO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_CMUX;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_CO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_CO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_DMUX;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_DO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_DO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_AO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_AO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_BO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_BO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_CO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_CO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_DO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_DO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D_XOR;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_A;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_A1;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_A2;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_A3;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_A4;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_A5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_A6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_AMUX;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_AO5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_AO6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_A_CY;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_A_XOR;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_B;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_B1;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_B2;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_B3;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_B4;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_B5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_B6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_BMUX;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_BO5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_BO6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_B_CY;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_B_XOR;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_C;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_C1;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_C2;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_C3;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_C4;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_C5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_C6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_CMUX;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_CO5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_CO6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_C_CY;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_C_XOR;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_D;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_D1;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_D2;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_D3;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_D4;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_D5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_D6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_DMUX;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_DO5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_DO6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_D_CY;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X0Y31_D_XOR;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_A;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_A1;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_A2;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_A3;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_A4;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_A5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_A6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_AO5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_AO6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_A_CY;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_A_XOR;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_B;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_B1;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_B2;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_B3;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_B4;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_B5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_B6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_BO5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_BO6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_B_CY;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_B_XOR;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_C;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_C1;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_C2;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_C3;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_C4;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_C5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_C6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_CO5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_CO6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_C_CY;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_C_XOR;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_D;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_D1;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_D2;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_D3;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_D4;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_D5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_D6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_DO5;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_DO6;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_D_CY;
  wire [0:0] CLBLL_L_X2Y31_SLICE_X1Y31_D_XOR;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE1;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S0;
  wire [0:0] CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S1;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_CE;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_I;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_CE;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_I;
  wire [0:0] CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y11_I;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y12_I;
  wire [0:0] LIOB33_X0Y13_IOB_X0Y13_I;
  wire [0:0] LIOB33_X0Y13_IOB_X0Y14_I;
  wire [0:0] LIOB33_X0Y15_IOB_X0Y15_I;
  wire [0:0] LIOB33_X0Y15_IOB_X0Y16_I;
  wire [0:0] LIOB33_X0Y17_IOB_X0Y17_I;
  wire [0:0] LIOB33_X0Y17_IOB_X0Y18_I;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y19_I;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y20_I;
  wire [0:0] LIOB33_X0Y21_IOB_X0Y21_I;
  wire [0:0] LIOB33_X0Y21_IOB_X0Y22_I;
  wire [0:0] LIOB33_X0Y23_IOB_X0Y23_I;
  wire [0:0] LIOB33_X0Y23_IOB_X0Y24_I;
  wire [0:0] LIOB33_X0Y25_IOB_X0Y25_I;
  wire [0:0] LIOB33_X0Y25_IOB_X0Y26_I;
  wire [0:0] LIOB33_X0Y27_IOB_X0Y27_I;
  wire [0:0] LIOB33_X0Y27_IOB_X0Y28_I;
  wire [0:0] LIOB33_X0Y29_IOB_X0Y29_I;
  wire [0:0] LIOB33_X0Y29_IOB_X0Y30_I;
  wire [0:0] LIOB33_X0Y31_IOB_X0Y31_I;
  wire [0:0] LIOB33_X0Y31_IOB_X0Y32_I;
  wire [0:0] LIOB33_X0Y33_IOB_X0Y33_I;
  wire [0:0] LIOB33_X0Y33_IOB_X0Y34_I;
  wire [0:0] LIOB33_X0Y35_IOB_X0Y35_I;
  wire [0:0] LIOB33_X0Y35_IOB_X0Y36_I;
  wire [0:0] LIOB33_X0Y37_IOB_X0Y37_I;
  wire [0:0] LIOB33_X0Y37_IOB_X0Y38_I;
  wire [0:0] LIOB33_X0Y39_IOB_X0Y39_I;
  wire [0:0] LIOB33_X0Y39_IOB_X0Y40_I;
  wire [0:0] LIOB33_X0Y41_IOB_X0Y41_I;
  wire [0:0] LIOB33_X0Y41_IOB_X0Y42_I;
  wire [0:0] LIOB33_X0Y43_IOB_X0Y43_I;
  wire [0:0] LIOB33_X0Y45_IOB_X0Y45_I;
  wire [0:0] LIOB33_X0Y45_IOB_X0Y46_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y10_I;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_CE1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_CLK;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_CLKB;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_Q1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_Q2;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_SR;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_CE1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_CLK;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_CLKB;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_Q1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_Q2;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_SR;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_CE1;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_CLK;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_CLKB;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_Q1;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_Q2;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_SR;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_CE1;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_CLK;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_CLKB;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_Q1;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_Q2;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_SR;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_CE1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_CLK;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_CLKB;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q2;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_SR;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_CE1;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_CLK;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_CLKB;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_Q1;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_Q2;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_SR;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_CE1;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_CLK;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_CLKB;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_Q1;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_Q2;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_SR;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_CE1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_CLK;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_CLKB;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q2;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_SR;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_CE1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_CLK;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_CLKB;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q2;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_SR;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_CE1;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_CLK;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_CLKB;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_Q1;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_Q2;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_SR;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_CE1;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_CLK;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_CLKB;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_Q1;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_Q2;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_SR;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y15_CE1;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y15_CLK;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y15_CLKB;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y15_D;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y15_Q1;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y15_Q2;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y15_SR;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y16_CE1;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y16_CLK;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y16_CLKB;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y16_D;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y16_Q1;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y16_Q2;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y16_SR;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y17_CE1;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y17_CLK;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y17_CLKB;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y17_D;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y17_Q1;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y17_Q2;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y17_SR;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y18_CE1;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y18_CLK;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y18_CLKB;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y18_D;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y18_Q1;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y18_Q2;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y18_SR;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y21_CE1;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y21_CLK;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y21_CLKB;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y21_D;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y21_Q1;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y21_Q2;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y21_SR;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y22_CE1;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y22_CLK;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y22_CLKB;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y22_D;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y22_Q1;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y22_Q2;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y22_SR;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y23_CE1;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y23_CLK;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y23_CLKB;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y23_D;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y23_Q1;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y23_Q2;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y23_SR;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y24_CE1;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y24_CLK;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y24_CLKB;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y24_D;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y24_Q1;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y24_Q2;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y24_SR;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y25_CE1;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y25_CLK;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y25_CLKB;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y25_D;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y25_Q1;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y25_Q2;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y25_SR;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y26_CE1;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y26_CLK;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y26_CLKB;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y26_D;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y26_Q1;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y26_Q2;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y26_SR;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y27_CE1;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y27_CLK;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y27_CLKB;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y27_D;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y27_Q1;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y27_Q2;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y27_SR;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y28_CE1;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y28_CLK;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y28_CLKB;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y28_D;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y28_Q1;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y28_Q2;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y28_SR;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y29_CE1;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y29_CLK;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y29_CLKB;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y29_D;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y29_Q1;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y29_Q2;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y29_SR;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y30_CE1;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y30_CLK;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y30_CLKB;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y30_D;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y30_Q1;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y30_Q2;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y30_SR;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y33_CE1;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y33_CLK;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y33_CLKB;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y33_D;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y33_Q1;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y33_Q2;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y33_SR;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y34_CE1;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y34_CLK;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y34_CLKB;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y34_D;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y34_Q1;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y34_Q2;
  wire [0:0] LIOI3_X0Y33_ILOGIC_X0Y34_SR;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y35_CE1;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y35_CLK;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y35_CLKB;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y35_D;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y35_Q1;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y35_Q2;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y35_SR;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y36_CE1;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y36_CLK;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y36_CLKB;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y36_D;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y36_Q1;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y36_Q2;
  wire [0:0] LIOI3_X0Y35_ILOGIC_X0Y36_SR;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y39_CE1;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y39_CLK;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y39_CLKB;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y39_D;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y39_Q1;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y39_Q2;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y39_SR;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y40_CE1;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y40_CLK;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y40_CLKB;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y40_D;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y40_Q1;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y40_Q2;
  wire [0:0] LIOI3_X0Y39_ILOGIC_X0Y40_SR;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y41_CE1;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y41_CLK;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y41_CLKB;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y41_D;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y41_Q1;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y41_Q2;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y41_SR;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y42_CE1;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y42_CLK;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y42_CLKB;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y42_D;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y42_Q1;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y42_Q2;
  wire [0:0] LIOI3_X0Y41_ILOGIC_X0Y42_SR;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y45_CE1;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y45_CLK;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y45_CLKB;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y45_D;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y45_Q1;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y45_Q2;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y45_SR;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y46_CE1;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y46_CLK;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y46_CLKB;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y46_D;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y46_Q1;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y46_Q2;
  wire [0:0] LIOI3_X0Y45_ILOGIC_X0Y46_SR;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_CE1;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_CLK;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_CLKB;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_Q1;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_Q2;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_SR;
  wire [0:0] RIOB33_X43Y23_IOB_X1Y24_I;
  wire [0:0] RIOB33_X43Y25_IOB_X1Y26_I;
  wire [0:0] RIOB33_X43Y43_IOB_X1Y43_O;
  wire [0:0] RIOB33_X43Y43_IOB_X1Y44_O;
  wire [0:0] RIOB33_X43Y45_IOB_X1Y45_I;
  wire [0:0] RIOB33_X43Y45_IOB_X1Y46_I;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_D1;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_OQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_T1;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_TQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_D1;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_OQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_T1;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_TQ;
  wire [0:0] RIOI3_X43Y23_ILOGIC_X1Y24_D;
  wire [0:0] RIOI3_X43Y23_ILOGIC_X1Y24_O;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_D;
  wire [0:0] RIOI3_X43Y25_ILOGIC_X1Y26_O;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y45_D;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y45_O;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y46_D;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y46_O;


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000101)
  ) CLBLL_L_X2Y22_SLICE_X0Y22_ALUT (
.I0(LIOI3_X0Y33_ILOGIC_X0Y34_Q2),
.I1(LIOI3_X0Y35_ILOGIC_X0Y36_Q2),
.I2(LIOI3_X0Y35_ILOGIC_X0Y35_Q2),
.I3(1'b1),
.I4(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q2),
.I5(1'b1),
.O5(CLBLL_L_X2Y22_SLICE_X0Y22_AO5),
.O6(CLBLL_L_X2Y22_SLICE_X0Y22_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000011)
  ) CLBLL_L_X2Y22_SLICE_X0Y22_BLUT (
.I0(LIOI3_X0Y35_ILOGIC_X0Y35_Q1),
.I1(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q1),
.I2(1'b1),
.I3(LIOI3_X0Y33_ILOGIC_X0Y34_Q1),
.I4(LIOI3_X0Y35_ILOGIC_X0Y36_Q1),
.I5(1'b1),
.O5(CLBLL_L_X2Y22_SLICE_X0Y22_BO5),
.O6(CLBLL_L_X2Y22_SLICE_X0Y22_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000000)
  ) CLBLL_L_X2Y22_SLICE_X0Y22_CLUT (
.I0(LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_Q2),
.I1(LIOI3_X0Y11_ILOGIC_X0Y12_Q2),
.I2(1'b1),
.I3(LIOI3_X0Y9_ILOGIC_X0Y10_Q2),
.I4(LIOI3_X0Y11_ILOGIC_X0Y11_Q2),
.I5(1'b1),
.O5(CLBLL_L_X2Y22_SLICE_X0Y22_CO5),
.O6(CLBLL_L_X2Y22_SLICE_X0Y22_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000000)
  ) CLBLL_L_X2Y22_SLICE_X0Y22_DLUT (
.I0(LIOI3_X0Y9_ILOGIC_X0Y10_Q1),
.I1(LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_Q1),
.I2(1'b1),
.I3(LIOI3_X0Y11_ILOGIC_X0Y12_Q1),
.I4(LIOI3_X0Y11_ILOGIC_X0Y11_Q1),
.I5(1'b1),
.O5(CLBLL_L_X2Y22_SLICE_X0Y22_DO5),
.O6(CLBLL_L_X2Y22_SLICE_X0Y22_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y22_SLICE_X1Y22_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y22_SLICE_X1Y22_AO5),
.O6(CLBLL_L_X2Y22_SLICE_X1Y22_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y22_SLICE_X1Y22_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y22_SLICE_X1Y22_BO5),
.O6(CLBLL_L_X2Y22_SLICE_X1Y22_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y22_SLICE_X1Y22_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y22_SLICE_X1Y22_CO5),
.O6(CLBLL_L_X2Y22_SLICE_X1Y22_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y22_SLICE_X1Y22_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y22_SLICE_X1Y22_DO5),
.O6(CLBLL_L_X2Y22_SLICE_X1Y22_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLL_L_X2Y24_SLICE_X0Y24_ALUT (
.I0(CLBLL_L_X2Y31_SLICE_X0Y31_CO6),
.I1(CLBLL_L_X2Y25_SLICE_X0Y25_CO6),
.I2(CLBLL_L_X2Y24_SLICE_X0Y24_DO6),
.I3(CLBLL_L_X2Y25_SLICE_X0Y25_AO5),
.I4(CLBLL_L_X2Y22_SLICE_X0Y22_AO5),
.I5(CLBLL_L_X2Y24_SLICE_X0Y24_BO6),
.O5(CLBLL_L_X2Y24_SLICE_X0Y24_AO5),
.O6(CLBLL_L_X2Y24_SLICE_X0Y24_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000000000000)
  ) CLBLL_L_X2Y24_SLICE_X0Y24_BLUT (
.I0(LIOI3_X0Y15_ILOGIC_X0Y15_Q2),
.I1(LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_Q2),
.I2(LIOI3_X0Y17_ILOGIC_X0Y17_Q2),
.I3(LIOI3_X0Y15_ILOGIC_X0Y16_Q2),
.I4(CLBLL_L_X2Y24_SLICE_X0Y24_CO6),
.I5(CLBLL_L_X2Y22_SLICE_X0Y22_CO6),
.O5(CLBLL_L_X2Y24_SLICE_X0Y24_BO5),
.O6(CLBLL_L_X2Y24_SLICE_X0Y24_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000500000000)
  ) CLBLL_L_X2Y24_SLICE_X0Y24_CLUT (
.I0(LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_Q2),
.I1(1'b1),
.I2(LIOI3_X0Y21_ILOGIC_X0Y21_Q2),
.I3(LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_Q2),
.I4(LIOI3_X0Y17_ILOGIC_X0Y18_Q2),
.I5(1'b1),
.O5(CLBLL_L_X2Y24_SLICE_X0Y24_CO5),
.O6(CLBLL_L_X2Y24_SLICE_X0Y24_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLL_L_X2Y24_SLICE_X0Y24_DLUT (
.I0(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q2),
.I1(LIOI3_X0Y39_ILOGIC_X0Y40_Q2),
.I2(LIOI3_X0Y39_ILOGIC_X0Y39_Q2),
.I3(CLBLL_L_X2Y31_SLICE_X0Y31_AO5),
.I4(LIOI3_X0Y41_ILOGIC_X0Y41_Q2),
.I5(1'b1),
.O5(CLBLL_L_X2Y24_SLICE_X0Y24_DO5),
.O6(CLBLL_L_X2Y24_SLICE_X0Y24_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h7fffffffffffffff)
  ) CLBLL_L_X2Y24_SLICE_X1Y24_ALUT (
.I0(CLBLL_L_X2Y31_SLICE_X0Y31_DO6),
.I1(CLBLL_L_X2Y25_SLICE_X0Y25_DO6),
.I2(CLBLL_L_X2Y24_SLICE_X1Y24_DO6),
.I3(CLBLL_L_X2Y25_SLICE_X0Y25_BO5),
.I4(CLBLL_L_X2Y22_SLICE_X0Y22_BO5),
.I5(CLBLL_L_X2Y24_SLICE_X1Y24_BO6),
.O5(CLBLL_L_X2Y24_SLICE_X1Y24_AO5),
.O6(CLBLL_L_X2Y24_SLICE_X1Y24_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0001000000000000)
  ) CLBLL_L_X2Y24_SLICE_X1Y24_BLUT (
.I0(LIOI3_X0Y15_ILOGIC_X0Y15_Q1),
.I1(LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_Q1),
.I2(LIOI3_X0Y17_ILOGIC_X0Y17_Q1),
.I3(LIOI3_X0Y15_ILOGIC_X0Y16_Q1),
.I4(CLBLL_L_X2Y24_SLICE_X1Y24_CO6),
.I5(CLBLL_L_X2Y22_SLICE_X0Y22_DO6),
.O5(CLBLL_L_X2Y24_SLICE_X1Y24_BO5),
.O6(CLBLL_L_X2Y24_SLICE_X1Y24_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000500000000)
  ) CLBLL_L_X2Y24_SLICE_X1Y24_CLUT (
.I0(LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_Q1),
.I1(1'b1),
.I2(LIOI3_X0Y21_ILOGIC_X0Y21_Q1),
.I3(LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_Q1),
.I4(LIOI3_X0Y17_ILOGIC_X0Y18_Q1),
.I5(1'b1),
.O5(CLBLL_L_X2Y24_SLICE_X1Y24_CO5),
.O6(CLBLL_L_X2Y24_SLICE_X1Y24_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000010000000000)
  ) CLBLL_L_X2Y24_SLICE_X1Y24_DLUT (
.I0(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q1),
.I1(LIOI3_X0Y39_ILOGIC_X0Y40_Q1),
.I2(LIOI3_X0Y39_ILOGIC_X0Y39_Q1),
.I3(CLBLL_L_X2Y31_SLICE_X0Y31_BO5),
.I4(LIOI3_X0Y41_ILOGIC_X0Y41_Q1),
.I5(1'b1),
.O5(CLBLL_L_X2Y24_SLICE_X1Y24_DO5),
.O6(CLBLL_L_X2Y24_SLICE_X1Y24_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000101)
  ) CLBLL_L_X2Y25_SLICE_X0Y25_ALUT (
.I0(LIOI3_X0Y29_ILOGIC_X0Y30_Q2),
.I1(LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_Q2),
.I2(LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_Q2),
.I3(1'b1),
.I4(LIOI3_X0Y33_ILOGIC_X0Y33_Q2),
.I5(1'b1),
.O5(CLBLL_L_X2Y25_SLICE_X0Y25_AO5),
.O6(CLBLL_L_X2Y25_SLICE_X0Y25_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000011)
  ) CLBLL_L_X2Y25_SLICE_X0Y25_BLUT (
.I0(LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_Q1),
.I1(LIOI3_X0Y33_ILOGIC_X0Y33_Q1),
.I2(1'b1),
.I3(LIOI3_X0Y29_ILOGIC_X0Y30_Q1),
.I4(LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_Q1),
.I5(1'b1),
.O5(CLBLL_L_X2Y25_SLICE_X0Y25_BO5),
.O6(CLBLL_L_X2Y25_SLICE_X0Y25_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000000)
  ) CLBLL_L_X2Y25_SLICE_X0Y25_CLUT (
.I0(LIOI3_X0Y25_ILOGIC_X0Y25_Q2),
.I1(LIOI3_X0Y23_ILOGIC_X0Y24_Q2),
.I2(1'b1),
.I3(LIOI3_X0Y21_ILOGIC_X0Y22_Q2),
.I4(LIOI3_X0Y23_ILOGIC_X0Y23_Q2),
.I5(1'b1),
.O5(CLBLL_L_X2Y25_SLICE_X0Y25_CO5),
.O6(CLBLL_L_X2Y25_SLICE_X0Y25_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000000)
  ) CLBLL_L_X2Y25_SLICE_X0Y25_DLUT (
.I0(LIOI3_X0Y21_ILOGIC_X0Y22_Q1),
.I1(LIOI3_X0Y25_ILOGIC_X0Y25_Q1),
.I2(1'b1),
.I3(LIOI3_X0Y23_ILOGIC_X0Y24_Q1),
.I4(LIOI3_X0Y23_ILOGIC_X0Y23_Q1),
.I5(1'b1),
.O5(CLBLL_L_X2Y25_SLICE_X0Y25_DO5),
.O6(CLBLL_L_X2Y25_SLICE_X0Y25_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y25_SLICE_X1Y25_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y25_SLICE_X1Y25_AO5),
.O6(CLBLL_L_X2Y25_SLICE_X1Y25_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y25_SLICE_X1Y25_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y25_SLICE_X1Y25_BO5),
.O6(CLBLL_L_X2Y25_SLICE_X1Y25_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y25_SLICE_X1Y25_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y25_SLICE_X1Y25_CO5),
.O6(CLBLL_L_X2Y25_SLICE_X1Y25_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y25_SLICE_X1Y25_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y25_SLICE_X1Y25_DO5),
.O6(CLBLL_L_X2Y25_SLICE_X1Y25_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000101)
  ) CLBLL_L_X2Y31_SLICE_X0Y31_ALUT (
.I0(LIOI3_X0Y41_ILOGIC_X0Y42_Q2),
.I1(LIOI3_X0Y45_ILOGIC_X0Y45_Q2),
.I2(LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q2),
.I3(1'b1),
.I4(LIOI3_X0Y45_ILOGIC_X0Y46_Q2),
.I5(1'b1),
.O5(CLBLL_L_X2Y31_SLICE_X0Y31_AO5),
.O6(CLBLL_L_X2Y31_SLICE_X0Y31_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000011)
  ) CLBLL_L_X2Y31_SLICE_X0Y31_BLUT (
.I0(LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q1),
.I1(LIOI3_X0Y45_ILOGIC_X0Y46_Q1),
.I2(1'b1),
.I3(LIOI3_X0Y41_ILOGIC_X0Y42_Q1),
.I4(LIOI3_X0Y45_ILOGIC_X0Y45_Q1),
.I5(1'b1),
.O5(CLBLL_L_X2Y31_SLICE_X0Y31_BO5),
.O6(CLBLL_L_X2Y31_SLICE_X0Y31_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000000)
  ) CLBLL_L_X2Y31_SLICE_X0Y31_CLUT (
.I0(LIOI3_X0Y29_ILOGIC_X0Y29_Q2),
.I1(LIOI3_X0Y27_ILOGIC_X0Y28_Q2),
.I2(1'b1),
.I3(LIOI3_X0Y25_ILOGIC_X0Y26_Q2),
.I4(LIOI3_X0Y27_ILOGIC_X0Y27_Q2),
.I5(1'b1),
.O5(CLBLL_L_X2Y31_SLICE_X0Y31_CO5),
.O6(CLBLL_L_X2Y31_SLICE_X0Y31_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000001100000000)
  ) CLBLL_L_X2Y31_SLICE_X0Y31_DLUT (
.I0(LIOI3_X0Y25_ILOGIC_X0Y26_Q1),
.I1(LIOI3_X0Y29_ILOGIC_X0Y29_Q1),
.I2(1'b1),
.I3(LIOI3_X0Y27_ILOGIC_X0Y28_Q1),
.I4(LIOI3_X0Y27_ILOGIC_X0Y27_Q1),
.I5(1'b1),
.O5(CLBLL_L_X2Y31_SLICE_X0Y31_DO5),
.O6(CLBLL_L_X2Y31_SLICE_X0Y31_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y31_SLICE_X1Y31_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y31_SLICE_X1Y31_AO5),
.O6(CLBLL_L_X2Y31_SLICE_X1Y31_AO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y31_SLICE_X1Y31_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y31_SLICE_X1Y31_BO5),
.O6(CLBLL_L_X2Y31_SLICE_X1Y31_BO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y31_SLICE_X1Y31_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y31_SLICE_X1Y31_CO5),
.O6(CLBLL_L_X2Y31_SLICE_X1Y31_CO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y31_SLICE_X1Y31_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y31_SLICE_X1Y31_DO5),
.O6(CLBLL_L_X2Y31_SLICE_X1Y31_DO6)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X43Y25_IOB_X1Y26_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFGCTRL" *)
  BUFGCTRL #(
    .INIT_OUT(0),
    .IS_CE0_INVERTED(0),
    .IS_CE1_INVERTED(1),
    .IS_IGNORE0_INVERTED(1),
    .IS_IGNORE1_INVERTED(0),
    .IS_S0_INVERTED(0),
    .IS_S1_INVERTED(1),
    .PRESELECT_I0("TRUE"),
    .PRESELECT_I1("FALSE")
  ) CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_BUFGCTRL (
.CE0(1'b1),
.CE1(1'b1),
.I0(RIOB33_X43Y23_IOB_X1Y24_I),
.I1(1'b1),
.IGNORE0(1'b1),
.IGNORE1(1'b1),
.O(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O),
.S0(1'b1),
.S1(1'b1)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O),
.O(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "BUFHCE" *)
  BUFHCE #(
    .CE_TYPE("SYNC"),
    .INIT_OUT(0),
    .IS_CE_INVERTED(0)
  ) CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_BUFHCE (
.CE(1'b1),
.I(CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O),
.O(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y9_IOB_X0Y10_IBUF (
.I(io[35]),
.O(LIOB33_X0Y9_IOB_X0Y10_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y11_IOB_X0Y11_IBUF (
.I(io[34]),
.O(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y11_IOB_X0Y12_IBUF (
.I(io[33]),
.O(LIOB33_X0Y11_IOB_X0Y12_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y13_IOB_X0Y13_IBUF (
.I(io[32]),
.O(LIOB33_X0Y13_IOB_X0Y13_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y13_IOB_X0Y14_IBUF (
.I(io[31]),
.O(LIOB33_X0Y13_IOB_X0Y14_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y15_IOB_X0Y15_IBUF (
.I(io[30]),
.O(LIOB33_X0Y15_IOB_X0Y15_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y15_IOB_X0Y16_IBUF (
.I(io[29]),
.O(LIOB33_X0Y15_IOB_X0Y16_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y17_IOB_X0Y17_IBUF (
.I(io[28]),
.O(LIOB33_X0Y17_IOB_X0Y17_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y17_IOB_X0Y18_IBUF (
.I(io[27]),
.O(LIOB33_X0Y17_IOB_X0Y18_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y19_IOB_X0Y19_IBUF (
.I(io[26]),
.O(LIOB33_X0Y19_IOB_X0Y19_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y19_IOB_X0Y20_IBUF (
.I(io[25]),
.O(LIOB33_X0Y19_IOB_X0Y20_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y21_IOB_X0Y21_IBUF (
.I(io[24]),
.O(LIOB33_X0Y21_IOB_X0Y21_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y21_IOB_X0Y22_IBUF (
.I(io[23]),
.O(LIOB33_X0Y21_IOB_X0Y22_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y23_IOB_X0Y23_IBUF (
.I(io[22]),
.O(LIOB33_X0Y23_IOB_X0Y23_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y23_IOB_X0Y24_IBUF (
.I(io[21]),
.O(LIOB33_X0Y23_IOB_X0Y24_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y25_IOB_X0Y25_IBUF (
.I(io[20]),
.O(LIOB33_X0Y25_IOB_X0Y25_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y25_IOB_X0Y26_IBUF (
.I(io[19]),
.O(LIOB33_X0Y25_IOB_X0Y26_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y27_IOB_X0Y27_IBUF (
.I(io[18]),
.O(LIOB33_X0Y27_IOB_X0Y27_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y27_IOB_X0Y28_IBUF (
.I(io[17]),
.O(LIOB33_X0Y27_IOB_X0Y28_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y29_IOB_X0Y29_IBUF (
.I(io[16]),
.O(LIOB33_X0Y29_IOB_X0Y29_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y29_IOB_X0Y30_IBUF (
.I(io[15]),
.O(LIOB33_X0Y29_IOB_X0Y30_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y31_IOB_X0Y31_IBUF (
.I(io[14]),
.O(LIOB33_X0Y31_IOB_X0Y31_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y31_IOB_X0Y32_IBUF (
.I(io[13]),
.O(LIOB33_X0Y31_IOB_X0Y32_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y33_IOB_X0Y33_IBUF (
.I(io[12]),
.O(LIOB33_X0Y33_IOB_X0Y33_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y33_IOB_X0Y34_IBUF (
.I(io[11]),
.O(LIOB33_X0Y33_IOB_X0Y34_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y35_IOB_X0Y35_IBUF (
.I(io[10]),
.O(LIOB33_X0Y35_IOB_X0Y35_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y35_IOB_X0Y36_IBUF (
.I(io[9]),
.O(LIOB33_X0Y35_IOB_X0Y36_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y37_IOB_X0Y37_IBUF (
.I(io[8]),
.O(LIOB33_X0Y37_IOB_X0Y37_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y37_IOB_X0Y38_IBUF (
.I(io[7]),
.O(LIOB33_X0Y37_IOB_X0Y38_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y39_IOB_X0Y39_IBUF (
.I(io[6]),
.O(LIOB33_X0Y39_IOB_X0Y39_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y39_IOB_X0Y40_IBUF (
.I(io[5]),
.O(LIOB33_X0Y39_IOB_X0Y40_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y41_IOB_X0Y41_IBUF (
.I(io[4]),
.O(LIOB33_X0Y41_IOB_X0Y41_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y41_IOB_X0Y42_IBUF (
.I(io[3]),
.O(LIOB33_X0Y41_IOB_X0Y42_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y43_IOB_X0Y43_IBUF (
.I(io[2]),
.O(LIOB33_X0Y43_IOB_X0Y43_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y45_IOB_X0Y45_IBUF (
.I(io[1]),
.O(LIOB33_X0Y45_IOB_X0Y45_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y45_IOB_X0Y46_IBUF (
.I(io[0]),
.O(LIOB33_X0Y45_IOB_X0Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y9_ILOGIC_X0Y10_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y9_IOB_X0Y10_I),
.Q1(LIOI3_X0Y9_ILOGIC_X0Y10_Q1),
.Q2(LIOI3_X0Y9_ILOGIC_X0Y10_Q2),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y11_ILOGIC_X0Y12_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y11_IOB_X0Y12_I),
.Q1(LIOI3_X0Y11_ILOGIC_X0Y12_Q1),
.Q2(LIOI3_X0Y11_ILOGIC_X0Y12_Q2),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y11_ILOGIC_X0Y11_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y11_IOB_X0Y11_I),
.Q1(LIOI3_X0Y11_ILOGIC_X0Y11_Q1),
.Q2(LIOI3_X0Y11_ILOGIC_X0Y11_Q2),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y15_ILOGIC_X0Y16_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y15_IOB_X0Y16_I),
.Q1(LIOI3_X0Y15_ILOGIC_X0Y16_Q1),
.Q2(LIOI3_X0Y15_ILOGIC_X0Y16_Q2),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y15_ILOGIC_X0Y15_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y15_IOB_X0Y15_I),
.Q1(LIOI3_X0Y15_ILOGIC_X0Y15_Q1),
.Q2(LIOI3_X0Y15_ILOGIC_X0Y15_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y17_ILOGIC_X0Y18_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y17_IOB_X0Y18_I),
.Q1(LIOI3_X0Y17_ILOGIC_X0Y18_Q1),
.Q2(LIOI3_X0Y17_ILOGIC_X0Y18_Q2),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y17_ILOGIC_X0Y17_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y17_IOB_X0Y17_I),
.Q1(LIOI3_X0Y17_ILOGIC_X0Y17_Q1),
.Q2(LIOI3_X0Y17_ILOGIC_X0Y17_Q2),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y21_ILOGIC_X0Y22_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y21_IOB_X0Y22_I),
.Q1(LIOI3_X0Y21_ILOGIC_X0Y22_Q1),
.Q2(LIOI3_X0Y21_ILOGIC_X0Y22_Q2),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y21_ILOGIC_X0Y21_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y21_IOB_X0Y21_I),
.Q1(LIOI3_X0Y21_ILOGIC_X0Y21_Q1),
.Q2(LIOI3_X0Y21_ILOGIC_X0Y21_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y23_ILOGIC_X0Y24_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y23_IOB_X0Y24_I),
.Q1(LIOI3_X0Y23_ILOGIC_X0Y24_Q1),
.Q2(LIOI3_X0Y23_ILOGIC_X0Y24_Q2),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y23_ILOGIC_X0Y23_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y23_IOB_X0Y23_I),
.Q1(LIOI3_X0Y23_ILOGIC_X0Y23_Q1),
.Q2(LIOI3_X0Y23_ILOGIC_X0Y23_Q2),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y25_ILOGIC_X0Y26_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y25_IOB_X0Y26_I),
.Q1(LIOI3_X0Y25_ILOGIC_X0Y26_Q1),
.Q2(LIOI3_X0Y25_ILOGIC_X0Y26_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y25_ILOGIC_X0Y25_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y25_IOB_X0Y25_I),
.Q1(LIOI3_X0Y25_ILOGIC_X0Y25_Q1),
.Q2(LIOI3_X0Y25_ILOGIC_X0Y25_Q2),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y27_ILOGIC_X0Y28_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y27_IOB_X0Y28_I),
.Q1(LIOI3_X0Y27_ILOGIC_X0Y28_Q1),
.Q2(LIOI3_X0Y27_ILOGIC_X0Y28_Q2),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_X0Y27_ILOGIC_X0Y27_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y27_IOB_X0Y27_I),
.Q1(LIOI3_X0Y27_ILOGIC_X0Y27_Q1),
.Q2(LIOI3_X0Y27_ILOGIC_X0Y27_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y29_ILOGIC_X0Y30_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y29_IOB_X0Y30_I),
.Q1(LIOI3_X0Y29_ILOGIC_X0Y30_Q1),
.Q2(LIOI3_X0Y29_ILOGIC_X0Y30_Q2),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y29_ILOGIC_X0Y29_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y29_IOB_X0Y29_I),
.Q1(LIOI3_X0Y29_ILOGIC_X0Y29_Q1),
.Q2(LIOI3_X0Y29_ILOGIC_X0Y29_Q2),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y33_ILOGIC_X0Y34_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y33_IOB_X0Y34_I),
.Q1(LIOI3_X0Y33_ILOGIC_X0Y34_Q1),
.Q2(LIOI3_X0Y33_ILOGIC_X0Y34_Q2),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y33_ILOGIC_X0Y33_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y33_IOB_X0Y33_I),
.Q1(LIOI3_X0Y33_ILOGIC_X0Y33_Q1),
.Q2(LIOI3_X0Y33_ILOGIC_X0Y33_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y35_ILOGIC_X0Y36_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y35_IOB_X0Y36_I),
.Q1(LIOI3_X0Y35_ILOGIC_X0Y36_Q1),
.Q2(LIOI3_X0Y35_ILOGIC_X0Y36_Q2),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y35_ILOGIC_X0Y35_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y35_IOB_X0Y35_I),
.Q1(LIOI3_X0Y35_ILOGIC_X0Y35_Q1),
.Q2(LIOI3_X0Y35_ILOGIC_X0Y35_Q2),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y39_ILOGIC_X0Y40_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y39_IOB_X0Y40_I),
.Q1(LIOI3_X0Y39_ILOGIC_X0Y40_Q1),
.Q2(LIOI3_X0Y39_ILOGIC_X0Y40_Q2),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y39_ILOGIC_X0Y39_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y39_IOB_X0Y39_I),
.Q1(LIOI3_X0Y39_ILOGIC_X0Y39_Q1),
.Q2(LIOI3_X0Y39_ILOGIC_X0Y39_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y41_ILOGIC_X0Y42_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y41_IOB_X0Y42_I),
.Q1(LIOI3_X0Y41_ILOGIC_X0Y42_Q1),
.Q2(LIOI3_X0Y41_ILOGIC_X0Y42_Q2),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y41_ILOGIC_X0Y41_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y41_IOB_X0Y41_I),
.Q1(LIOI3_X0Y41_ILOGIC_X0Y41_Q1),
.Q2(LIOI3_X0Y41_ILOGIC_X0Y41_Q2),
.S(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y45_ILOGIC_X0Y46_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y45_IOB_X0Y46_I),
.Q1(LIOI3_X0Y45_ILOGIC_X0Y46_Q1),
.Q2(LIOI3_X0Y45_ILOGIC_X0Y46_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_X0Y45_ILOGIC_X0Y45_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y45_IOB_X0Y45_I),
.Q1(LIOI3_X0Y45_ILOGIC_X0Y45_Q1),
.Q2(LIOI3_X0Y45_ILOGIC_X0Y45_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y19_IOB_X0Y20_I),
.Q1(LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_Q1),
.Q2(LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y19_IOB_X0Y19_I),
.Q1(LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_Q1),
.Q2(LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_Q2),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y31_IOB_X0Y32_I),
.Q1(LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_Q1),
.Q2(LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y31_IOB_X0Y31_I),
.Q1(LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_Q1),
.Q2(LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_Q2),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y43_IOB_X0Y43_I),
.Q1(LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q1),
.Q2(LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q2),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y13_IOB_X0Y14_I),
.Q1(LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_Q1),
.Q2(LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("OPPOSITE_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("SYNC")
  ) LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y13_IOB_X0Y13_I),
.Q1(LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_Q1),
.Q2(LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_Q2),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b1),
    .INIT_Q2(1'b0),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y37_IOB_X0Y38_I),
.Q1(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q1),
.Q2(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q2),
.R(1'b0),
.S(1'b0)
  );


  (* KEEP, DONT_TOUCH, BEL = "IFF" *)
  IDDR_2CLK #(
    .DDR_CLK_EDGE("SAME_EDGE"),
    .INIT_Q1(1'b0),
    .INIT_Q2(1'b1),
    .IS_C_INVERTED(1'b0),
    .IS_D_INVERTED(1'b0),
    .SRTYPE("ASYNC")
  ) LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_IDDR_2CLK (
.C(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O),
.CB(CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O),
.CE(RIOB33_X43Y45_IOB_X1Y45_I),
.D(LIOB33_X0Y37_IOB_X0Y37_I),
.Q1(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q1),
.Q2(LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q2),
.R(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y23_IOB_X1Y24_IBUF (
.I(i_clkb),
.O(RIOB33_X43Y23_IOB_X1Y24_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y25_IOB_X1Y26_IBUF (
.I(i_clk),
.O(RIOB33_X43Y25_IOB_X1Y26_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y43_IOB_X1Y43_OBUF (
.I(CLBLL_L_X2Y24_SLICE_X0Y24_AO6),
.O(o_q2)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y43_IOB_X1Y44_OBUF (
.I(CLBLL_L_X2Y24_SLICE_X1Y24_AO6),
.O(o_q1)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y45_IOB_X1Y45_IBUF (
.I(i_ce),
.O(RIOB33_X43Y45_IOB_X1Y45_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y45_IOB_X1Y46_IBUF (
.I(i_rst),
.O(RIOB33_X43Y45_IOB_X1Y46_I)
  );
  assign CLBLL_L_X2Y22_SLICE_X0Y22_A = CLBLL_L_X2Y22_SLICE_X0Y22_AO6;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_B = CLBLL_L_X2Y22_SLICE_X0Y22_BO6;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_C = CLBLL_L_X2Y22_SLICE_X0Y22_CO6;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_D = CLBLL_L_X2Y22_SLICE_X0Y22_DO6;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_AMUX = CLBLL_L_X2Y22_SLICE_X0Y22_AO5;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_BMUX = CLBLL_L_X2Y22_SLICE_X0Y22_BO5;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_CMUX = CLBLL_L_X2Y22_SLICE_X0Y22_CO6;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_DMUX = CLBLL_L_X2Y22_SLICE_X0Y22_DO6;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_A = CLBLL_L_X2Y22_SLICE_X1Y22_AO6;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_B = CLBLL_L_X2Y22_SLICE_X1Y22_BO6;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_C = CLBLL_L_X2Y22_SLICE_X1Y22_CO6;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_D = CLBLL_L_X2Y22_SLICE_X1Y22_DO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_A = CLBLL_L_X2Y24_SLICE_X0Y24_AO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_B = CLBLL_L_X2Y24_SLICE_X0Y24_BO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_C = CLBLL_L_X2Y24_SLICE_X0Y24_CO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_D = CLBLL_L_X2Y24_SLICE_X0Y24_DO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_AMUX = CLBLL_L_X2Y24_SLICE_X0Y24_AO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_BMUX = CLBLL_L_X2Y24_SLICE_X0Y24_BO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_CMUX = CLBLL_L_X2Y24_SLICE_X0Y24_CO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_DMUX = CLBLL_L_X2Y24_SLICE_X0Y24_DO6;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_A = CLBLL_L_X2Y24_SLICE_X1Y24_AO6;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_B = CLBLL_L_X2Y24_SLICE_X1Y24_BO6;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_C = CLBLL_L_X2Y24_SLICE_X1Y24_CO6;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_D = CLBLL_L_X2Y24_SLICE_X1Y24_DO6;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_AMUX = CLBLL_L_X2Y24_SLICE_X1Y24_AO6;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_BMUX = CLBLL_L_X2Y24_SLICE_X1Y24_BO6;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_CMUX = CLBLL_L_X2Y24_SLICE_X1Y24_CO6;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_DMUX = CLBLL_L_X2Y24_SLICE_X1Y24_DO6;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_A = CLBLL_L_X2Y25_SLICE_X0Y25_AO6;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_B = CLBLL_L_X2Y25_SLICE_X0Y25_BO6;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_C = CLBLL_L_X2Y25_SLICE_X0Y25_CO6;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_D = CLBLL_L_X2Y25_SLICE_X0Y25_DO6;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_AMUX = CLBLL_L_X2Y25_SLICE_X0Y25_AO5;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_BMUX = CLBLL_L_X2Y25_SLICE_X0Y25_BO5;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_CMUX = CLBLL_L_X2Y25_SLICE_X0Y25_CO6;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_DMUX = CLBLL_L_X2Y25_SLICE_X0Y25_DO6;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_A = CLBLL_L_X2Y25_SLICE_X1Y25_AO6;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_B = CLBLL_L_X2Y25_SLICE_X1Y25_BO6;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_C = CLBLL_L_X2Y25_SLICE_X1Y25_CO6;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_D = CLBLL_L_X2Y25_SLICE_X1Y25_DO6;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_A = CLBLL_L_X2Y31_SLICE_X0Y31_AO6;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_B = CLBLL_L_X2Y31_SLICE_X0Y31_BO6;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_C = CLBLL_L_X2Y31_SLICE_X0Y31_CO6;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_D = CLBLL_L_X2Y31_SLICE_X0Y31_DO6;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_AMUX = CLBLL_L_X2Y31_SLICE_X0Y31_AO5;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_BMUX = CLBLL_L_X2Y31_SLICE_X0Y31_BO5;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_CMUX = CLBLL_L_X2Y31_SLICE_X0Y31_CO6;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_DMUX = CLBLL_L_X2Y31_SLICE_X0Y31_DO6;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_A = CLBLL_L_X2Y31_SLICE_X1Y31_AO6;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_B = CLBLL_L_X2Y31_SLICE_X1Y31_BO6;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_C = CLBLL_L_X2Y31_SLICE_X1Y31_CO6;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_D = CLBLL_L_X2Y31_SLICE_X1Y31_DO6;
  assign RIOI3_X43Y23_ILOGIC_X1Y24_O = RIOI3_X43Y23_ILOGIC_X1Y24_D;
  assign RIOI3_X43Y25_ILOGIC_X1Y26_O = RIOI3_X43Y25_ILOGIC_X1Y26_D;
  assign RIOI3_X43Y45_ILOGIC_X1Y46_O = RIOI3_X43Y45_ILOGIC_X1Y46_D;
  assign RIOI3_X43Y45_ILOGIC_X1Y45_O = RIOI3_X43Y45_ILOGIC_X1Y45_D;
  assign RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_OQ = RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_D1;
  assign RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_TQ = RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y44_T1;
  assign RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_OQ = RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_D1;
  assign RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_TQ = RIOI3_TBYTESRC_X43Y43_OLOGIC_X1Y43_T1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_C4 = LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_Q1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_C5 = LIOI3_X0Y17_ILOGIC_X0Y18_Q1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_C6 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y39_ILOGIC_X0Y40_D = LIOB33_X0Y39_IOB_X0Y40_I;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_D1 = LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_D2 = LIOI3_X0Y39_ILOGIC_X0Y40_Q1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_D3 = LIOI3_X0Y39_ILOGIC_X0Y39_Q1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_D4 = CLBLL_L_X2Y31_SLICE_X0Y31_BO5;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_D5 = LIOI3_X0Y41_ILOGIC_X0Y41_Q1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_D6 = 1'b1;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_D = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y39_ILOGIC_X0Y39_D = LIOB33_X0Y39_IOB_X0Y39_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_A1 = LIOI3_X0Y41_ILOGIC_X0Y42_Q2;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_A2 = LIOI3_X0Y45_ILOGIC_X0Y45_Q2;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_A3 = LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q2;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_A4 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_A5 = LIOI3_X0Y45_ILOGIC_X0Y46_Q2;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_A6 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_B1 = LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_Q1;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_B2 = LIOI3_X0Y45_ILOGIC_X0Y46_Q1;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_B3 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_B4 = LIOI3_X0Y41_ILOGIC_X0Y42_Q1;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_B5 = LIOI3_X0Y45_ILOGIC_X0Y45_Q1;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_B6 = 1'b1;
  assign LIOI3_X0Y33_ILOGIC_X0Y34_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y33_ILOGIC_X0Y34_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y33_ILOGIC_X0Y34_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_C1 = LIOI3_X0Y29_ILOGIC_X0Y29_Q2;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_C2 = LIOI3_X0Y27_ILOGIC_X0Y28_Q2;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_C3 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_C4 = LIOI3_X0Y25_ILOGIC_X0Y26_Q2;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_C5 = LIOI3_X0Y27_ILOGIC_X0Y27_Q2;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_C6 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_C3 = LIOI3_X0Y21_ILOGIC_X0Y21_Q1;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_D1 = LIOI3_X0Y25_ILOGIC_X0Y26_Q1;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_D2 = LIOI3_X0Y29_ILOGIC_X0Y29_Q1;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_D3 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_D4 = LIOI3_X0Y27_ILOGIC_X0Y28_Q1;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_D5 = LIOI3_X0Y27_ILOGIC_X0Y27_Q1;
  assign CLBLL_L_X2Y31_SLICE_X0Y31_D6 = 1'b1;
  assign LIOI3_X0Y33_ILOGIC_X0Y34_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y33_ILOGIC_X0Y33_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y33_ILOGIC_X0Y33_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y33_ILOGIC_X0Y33_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y33_ILOGIC_X0Y33_SR = 1'b0;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_A1 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_A2 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_A3 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_A4 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_A5 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_A6 = 1'b1;
  assign LIOI3_X0Y27_ILOGIC_X0Y28_D = LIOB33_X0Y27_IOB_X0Y28_I;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_B1 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_B2 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_B3 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_B4 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_B5 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_B6 = 1'b1;
  assign LIOI3_X0Y27_ILOGIC_X0Y27_D = LIOB33_X0Y27_IOB_X0Y27_I;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_C1 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_C2 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_C3 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_C4 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_C5 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_C6 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_D1 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_D2 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_D3 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_D4 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_D5 = 1'b1;
  assign CLBLL_L_X2Y31_SLICE_X1Y31_D6 = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_O;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_I = CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_O;
  assign LIOI3_X0Y23_ILOGIC_X0Y24_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y23_ILOGIC_X0Y24_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y23_ILOGIC_X0Y24_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y23_ILOGIC_X0Y24_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y23_ILOGIC_X0Y23_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y23_ILOGIC_X0Y23_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y23_ILOGIC_X0Y23_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y23_ILOGIC_X0Y23_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y17_ILOGIC_X0Y18_D = LIOB33_X0Y17_IOB_X0Y18_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE1 = 1'b1;
  assign LIOI3_X0Y17_ILOGIC_X0Y17_D = LIOB33_X0Y17_IOB_X0Y17_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S0 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_D = LIOB33_X0Y37_IOB_X0Y38_I;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_D = LIOB33_X0Y37_IOB_X0Y37_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_S1 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_A1 = LIOI3_X0Y29_ILOGIC_X0Y30_Q2;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_A2 = LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_Q2;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_A3 = LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_Q2;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_A4 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_A5 = LIOI3_X0Y33_ILOGIC_X0Y33_Q2;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_D = LIOB33_X0Y31_IOB_X0Y32_I;
  assign LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_D = LIOB33_X0Y31_IOB_X0Y31_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_B1 = LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_Q1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_B2 = LIOI3_X0Y33_ILOGIC_X0Y33_Q1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_B3 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_B4 = LIOI3_X0Y29_ILOGIC_X0Y30_Q1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_B5 = LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_Q1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_B6 = 1'b1;
  assign LIOI3_X0Y41_ILOGIC_X0Y42_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y41_ILOGIC_X0Y42_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_C1 = LIOI3_X0Y25_ILOGIC_X0Y25_Q2;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_C2 = LIOI3_X0Y23_ILOGIC_X0Y24_Q2;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_C3 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_C4 = LIOI3_X0Y21_ILOGIC_X0Y22_Q2;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_C5 = LIOI3_X0Y23_ILOGIC_X0Y23_Q2;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_C6 = 1'b1;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y41_ILOGIC_X0Y42_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y41_ILOGIC_X0Y41_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_D1 = LIOI3_X0Y21_ILOGIC_X0Y22_Q1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_D2 = LIOI3_X0Y25_ILOGIC_X0Y25_Q1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_D3 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_D4 = LIOI3_X0Y23_ILOGIC_X0Y24_Q1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_D5 = LIOI3_X0Y23_ILOGIC_X0Y23_Q1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_D6 = 1'b1;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y41_ILOGIC_X0Y41_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y45_ILOGIC_X0Y45_SR = 1'b0;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_A1 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_A2 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_A3 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_A4 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_A5 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_A6 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_IGNORE0 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_B1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_CE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_IGNORE1 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S0 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_S1 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_B2 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_B3 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_B4 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_B5 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_B6 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_C1 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_C2 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_C3 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_C4 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_A1 = LIOI3_X0Y33_ILOGIC_X0Y34_Q2;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_A2 = LIOI3_X0Y35_ILOGIC_X0Y36_Q2;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_A3 = LIOI3_X0Y35_ILOGIC_X0Y35_Q2;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_A4 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_A5 = LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q2;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_A6 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_C5 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_C6 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_B1 = LIOI3_X0Y35_ILOGIC_X0Y35_Q1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_D4 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_D5 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_D6 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_B2 = LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_Q1;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_B3 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_B4 = LIOI3_X0Y33_ILOGIC_X0Y34_Q1;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_B5 = LIOI3_X0Y35_ILOGIC_X0Y36_Q1;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_B6 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_C1 = LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_Q2;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_C2 = LIOI3_X0Y11_ILOGIC_X0Y12_Q2;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_C3 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_C4 = LIOI3_X0Y9_ILOGIC_X0Y10_Q2;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_C5 = LIOI3_X0Y11_ILOGIC_X0Y11_Q2;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_C6 = 1'b1;
  assign LIOI3_X0Y29_ILOGIC_X0Y30_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_D1 = LIOI3_X0Y9_ILOGIC_X0Y10_Q1;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_D2 = LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_Q1;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_D3 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_D4 = LIOI3_X0Y11_ILOGIC_X0Y12_Q1;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_D5 = LIOI3_X0Y11_ILOGIC_X0Y11_Q1;
  assign CLBLL_L_X2Y22_SLICE_X0Y22_D6 = 1'b1;
  assign LIOI3_X0Y29_ILOGIC_X0Y29_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y29_ILOGIC_X0Y29_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y29_ILOGIC_X0Y29_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_D = LIOB33_X0Y43_IOB_X0Y43_I;
  assign LIOI3_X0Y29_ILOGIC_X0Y29_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_A1 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_A2 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_A3 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_A4 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_A5 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_A6 = 1'b1;
  assign LIOI3_X0Y25_ILOGIC_X0Y26_D = LIOB33_X0Y25_IOB_X0Y26_I;
  assign LIOI3_X0Y25_ILOGIC_X0Y25_D = LIOB33_X0Y25_IOB_X0Y25_I;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_B1 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_B2 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_B3 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_B4 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_B5 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_B6 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_C1 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_C2 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_C3 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_C4 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_C5 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_C6 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_D1 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_D2 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_D3 = 1'b1;
  assign LIOI3_X0Y21_ILOGIC_X0Y22_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_D4 = 1'b1;
  assign LIOI3_X0Y21_ILOGIC_X0Y22_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y21_ILOGIC_X0Y22_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_D5 = 1'b1;
  assign CLBLL_L_X2Y22_SLICE_X1Y22_D6 = 1'b1;
  assign LIOI3_X0Y41_ILOGIC_X0Y42_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y21_ILOGIC_X0Y22_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y21_ILOGIC_X0Y21_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y21_ILOGIC_X0Y21_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y21_ILOGIC_X0Y21_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y21_ILOGIC_X0Y21_SR = 1'b0;
  assign LIOI3_X0Y45_ILOGIC_X0Y46_D = LIOB33_X0Y45_IOB_X0Y46_I;
  assign LIOI3_X0Y45_ILOGIC_X0Y45_D = LIOB33_X0Y45_IOB_X0Y45_I;
  assign LIOI3_TBYTESRC_X0Y43_ILOGIC_X0Y43_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign RIOB33_X43Y43_IOB_X1Y43_O = CLBLL_L_X2Y24_SLICE_X0Y24_AO6;
  assign RIOB33_X43Y43_IOB_X1Y44_O = CLBLL_L_X2Y24_SLICE_X1Y24_AO6;
  assign LIOI3_X0Y15_ILOGIC_X0Y16_D = LIOB33_X0Y15_IOB_X0Y16_I;
  assign LIOI3_X0Y15_ILOGIC_X0Y15_D = LIOB33_X0Y15_IOB_X0Y15_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_D = LIOB33_X0Y13_IOB_X0Y14_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_D = LIOB33_X0Y13_IOB_X0Y13_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_D = LIOB33_X0Y19_IOB_X0Y20_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_D = LIOB33_X0Y19_IOB_X0Y19_I;
  assign LIOI3_X0Y39_ILOGIC_X0Y40_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y39_ILOGIC_X0Y40_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y39_ILOGIC_X0Y40_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y39_ILOGIC_X0Y40_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y39_ILOGIC_X0Y39_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y39_ILOGIC_X0Y39_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y39_ILOGIC_X0Y39_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y41_ILOGIC_X0Y41_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y41_ILOGIC_X0Y41_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_SR = 1'b0;
  assign LIOI3_X0Y39_ILOGIC_X0Y39_SR = 1'b0;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y33_ILOGIC_X0Y34_D = LIOB33_X0Y33_IOB_X0Y34_I;
  assign LIOI3_X0Y33_ILOGIC_X0Y33_D = LIOB33_X0Y33_IOB_X0Y33_I;
  assign LIOI3_X0Y27_ILOGIC_X0Y28_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y27_ILOGIC_X0Y28_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y27_ILOGIC_X0Y28_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y27_ILOGIC_X0Y28_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y27_ILOGIC_X0Y27_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y27_ILOGIC_X0Y27_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y27_ILOGIC_X0Y27_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y27_ILOGIC_X0Y27_SR = 1'b0;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_D1 = 1'b1;
  assign LIOI3_X0Y23_ILOGIC_X0Y24_D = LIOB33_X0Y23_IOB_X0Y24_I;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_D2 = 1'b1;
  assign LIOI3_X0Y23_ILOGIC_X0Y23_D = LIOB33_X0Y23_IOB_X0Y23_I;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_D3 = 1'b1;
  assign LIOI3_X0Y35_ILOGIC_X0Y36_D = LIOB33_X0Y35_IOB_X0Y36_I;
  assign LIOI3_X0Y17_ILOGIC_X0Y18_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y17_ILOGIC_X0Y18_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y17_ILOGIC_X0Y18_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y35_ILOGIC_X0Y35_D = LIOB33_X0Y35_IOB_X0Y35_I;
  assign LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y17_ILOGIC_X0Y18_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y17_ILOGIC_X0Y17_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y17_ILOGIC_X0Y17_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y17_ILOGIC_X0Y17_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_SR = 1'b0;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y32_SR = 1'b0;
  assign LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y17_ILOGIC_X0Y17_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y37_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y41_ILOGIC_X0Y42_D = LIOB33_X0Y41_IOB_X0Y42_I;
  assign LIOI3_X0Y41_ILOGIC_X0Y41_D = LIOB33_X0Y41_IOB_X0Y41_I;
  assign LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_D = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_D = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y35_ILOGIC_X0Y36_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y35_ILOGIC_X0Y36_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_CE = 1'b1;
  assign CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_CE = 1'b1;
  assign LIOI3_X0Y35_ILOGIC_X0Y36_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y29_ILOGIC_X0Y30_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y29_ILOGIC_X0Y30_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y35_ILOGIC_X0Y36_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y29_ILOGIC_X0Y30_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y35_ILOGIC_X0Y35_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y35_ILOGIC_X0Y35_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y35_ILOGIC_X0Y35_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y35_ILOGIC_X0Y35_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_X0Y29_ILOGIC_X0Y30_D = LIOB33_X0Y29_IOB_X0Y30_I;
  assign LIOI3_X0Y29_ILOGIC_X0Y29_D = LIOB33_X0Y29_IOB_X0Y29_I;
  assign LIOI3_X0Y25_ILOGIC_X0Y26_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y25_ILOGIC_X0Y26_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y25_ILOGIC_X0Y26_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y25_ILOGIC_X0Y26_SR = 1'b0;
  assign LIOI3_X0Y25_ILOGIC_X0Y25_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y25_ILOGIC_X0Y25_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y25_ILOGIC_X0Y25_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y25_ILOGIC_X0Y25_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_A1 = CLBLL_L_X2Y31_SLICE_X0Y31_CO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_A2 = CLBLL_L_X2Y25_SLICE_X0Y25_CO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_A3 = CLBLL_L_X2Y24_SLICE_X0Y24_DO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_A4 = CLBLL_L_X2Y25_SLICE_X0Y25_AO5;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_A5 = CLBLL_L_X2Y22_SLICE_X0Y22_AO5;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_A6 = CLBLL_L_X2Y24_SLICE_X0Y24_BO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_B1 = LIOI3_X0Y15_ILOGIC_X0Y15_Q2;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_B2 = LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_Q2;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_B3 = LIOI3_X0Y17_ILOGIC_X0Y17_Q2;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_B4 = LIOI3_X0Y15_ILOGIC_X0Y16_Q2;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_B5 = CLBLL_L_X2Y24_SLICE_X0Y24_CO6;
  assign LIOI3_X0Y21_ILOGIC_X0Y22_D = LIOB33_X0Y21_IOB_X0Y22_I;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_B6 = CLBLL_L_X2Y22_SLICE_X0Y22_CO6;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I0 = RIOB33_X43Y25_IOB_X1Y26_I;
  assign LIOI3_X0Y21_ILOGIC_X0Y21_D = LIOB33_X0Y21_IOB_X0Y21_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y0_I1 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_C1 = LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_Q2;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_C2 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_C3 = LIOI3_X0Y21_ILOGIC_X0Y21_Q2;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_C4 = LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_Q2;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_C5 = LIOI3_X0Y17_ILOGIC_X0Y18_Q2;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_C6 = 1'b1;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I0 = RIOB33_X43Y23_IOB_X1Y24_I;
  assign CLK_BUFG_BOT_R_X60Y48_BUFGCTRL_X0Y1_I1 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_D1 = LIOI3_TBYTETERM_X0Y37_ILOGIC_X0Y38_Q2;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_D2 = LIOI3_X0Y39_ILOGIC_X0Y40_Q2;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_D3 = LIOI3_X0Y39_ILOGIC_X0Y39_Q2;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_D4 = CLBLL_L_X2Y31_SLICE_X0Y31_AO5;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_D5 = LIOI3_X0Y41_ILOGIC_X0Y41_Q2;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_D6 = 1'b1;
  assign LIOI3_X0Y45_ILOGIC_X0Y46_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y45_ILOGIC_X0Y46_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y45_ILOGIC_X0Y46_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y15_ILOGIC_X0Y16_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y15_ILOGIC_X0Y16_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y15_ILOGIC_X0Y16_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y45_ILOGIC_X0Y46_SR = 1'b0;
  assign LIOI3_X0Y45_ILOGIC_X0Y45_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y45_ILOGIC_X0Y45_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y45_ILOGIC_X0Y45_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign LIOI3_X0Y15_ILOGIC_X0Y16_SR = RIOB33_X43Y45_IOB_X1Y46_I;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_A1 = CLBLL_L_X2Y31_SLICE_X0Y31_DO6;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_A2 = CLBLL_L_X2Y25_SLICE_X0Y25_DO6;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_A3 = CLBLL_L_X2Y24_SLICE_X1Y24_DO6;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_A4 = CLBLL_L_X2Y25_SLICE_X0Y25_BO5;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_A5 = CLBLL_L_X2Y22_SLICE_X0Y22_BO5;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_A6 = CLBLL_L_X2Y24_SLICE_X1Y24_BO6;
  assign LIOI3_X0Y15_ILOGIC_X0Y15_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_X0Y15_ILOGIC_X0Y15_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign LIOI3_X0Y15_ILOGIC_X0Y15_CLKB = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y8_O;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_B1 = LIOI3_X0Y15_ILOGIC_X0Y15_Q1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_B2 = LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_Q1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_B3 = LIOI3_X0Y17_ILOGIC_X0Y17_Q1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_B4 = LIOI3_X0Y15_ILOGIC_X0Y16_Q1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_B5 = CLBLL_L_X2Y24_SLICE_X1Y24_CO6;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_B6 = CLBLL_L_X2Y22_SLICE_X0Y22_DO6;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_SR = 1'b0;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_CE1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_CLK = CLK_HROW_BOT_R_X60Y26_BUFHCE_X0Y9_O;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_C1 = LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_Q1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_C2 = 1'b1;
  assign LIOI3_X0Y15_ILOGIC_X0Y15_SR = 1'b0;
endmodule
