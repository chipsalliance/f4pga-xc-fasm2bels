// Copyright (C) 2021  The SymbiFlow Authors.
//
// Use of this source code is governed by a ISC-style
// license that can be found in the LICENSE file or at
// https://opensource.org/licenses/ISC
//
// SPDX-License-Identifier: ISC

module top(
  input rx,
  input [15:0] sw,
  output [15:0] led,
  output tx
  );
  wire [0:0] LIOB33_SING_X0Y0_IOB_X0Y0_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y111_O;
  wire [0:0] LIOB33_X0Y111_IOB_X0Y112_I;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y11_I;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y12_I;
  wire [0:0] LIOB33_X0Y17_IOB_X0Y18_O;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y19_O;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y20_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_O;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y2_O;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y3_O;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y4_O;
  wire [0:0] LIOB33_X0Y43_IOB_X0Y43_O;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y5_I;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y6_I;
  wire [0:0] LIOB33_X0Y7_IOB_X0Y7_I;
  wire [0:0] LIOB33_X0Y7_IOB_X0Y8_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y10_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y9_I;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_D1;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_OQ;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_T1;
  wire [0:0] LIOI3_SING_X0Y0_OLOGIC_X0Y0_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_O;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_D;
  wire [0:0] LIOI3_X0Y111_ILOGIC_X0Y112_O;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_D1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_OQ;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_T1;
  wire [0:0] LIOI3_X0Y111_OLOGIC_X0Y111_TQ;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_O;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_O;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_D1;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_OQ;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_T1;
  wire [0:0] LIOI3_X0Y17_OLOGIC_X0Y18_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y1_TQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_D1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_OQ;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_T1;
  wire [0:0] LIOI3_X0Y1_OLOGIC_X0Y2_TQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_D1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_OQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_T1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y3_TQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_D1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_OQ;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_T1;
  wire [0:0] LIOI3_X0Y3_OLOGIC_X0Y4_TQ;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y5_D;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y5_O;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_D;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_O;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_O;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y9_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y9_O;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERECRCCHECKEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERECRCGENEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERINTERRUPTMSGNUM0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERINTERRUPTMSGNUM1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERINTERRUPTMSGNUM2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERINTERRUPTMSGNUM3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERINTERRUPTMSGNUM4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERROOTERRCORRERRRECEIVED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERROOTERRCORRERRREPORTINGEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERROOTERRFATALERRRECEIVED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERROOTERRFATALERRREPORTINGEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERROOTERRNONFATALERRRECEIVED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERROOTERRNONFATALERRREPORTINGEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGBRIDGESERREN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGCOMMANDBUSMASTERENABLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGCOMMANDINTERRUPTDISABLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGCOMMANDIOENABLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGCOMMANDMEMENABLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGCOMMANDSERREN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2ARIFORWARDEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2ATOMICEGRESSBLOCK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2ATOMICREQUESTEREN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2CPLTIMEOUTDIS;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2CPLTIMEOUTVAL0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2CPLTIMEOUTVAL1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2CPLTIMEOUTVAL2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2CPLTIMEOUTVAL3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2IDOCPLEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2IDOREQEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2LTREN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2TLPPREFIXBLOCK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLAUXPOWEREN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLCORRERRREPORTINGEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLENABLERO;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLEXTTAGEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLFATALERRREPORTINGEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLMAXPAYLOAD0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLMAXPAYLOAD1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLMAXPAYLOAD2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLMAXREADREQ0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLMAXREADREQ1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLMAXREADREQ2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLNONFATALREPORTINGEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLNOSNOOPEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLPHANTOMEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLURERRREPORTINGEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVSTATUSCORRERRDETECTED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVSTATUSFATALERRDETECTED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVSTATUSNONFATALERRDETECTED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVSTATUSURDETECTED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSDEVICENUMBER0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSDEVICENUMBER1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSDEVICENUMBER2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSDEVICENUMBER3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSDEVICENUMBER4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSFUNCTIONNUMBER0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSFUNCTIONNUMBER1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSFUNCTIONNUMBER2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN32;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN33;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN34;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN35;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN36;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN37;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN38;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN39;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN40;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN41;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN42;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN43;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN44;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN45;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN46;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN47;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN48;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN49;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN50;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN51;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN52;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN53;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN54;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN55;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN56;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN57;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN58;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN59;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN60;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN61;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN62;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN63;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRACSN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG100;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG101;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG102;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG103;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG104;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG105;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG106;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG107;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG108;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG109;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG110;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG111;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG112;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG113;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG114;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG115;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG116;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG117;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG118;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG119;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG120;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG121;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG122;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG123;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG124;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG125;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG126;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG127;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG32;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG33;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG34;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG35;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG36;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG37;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG38;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG39;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG40;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG41;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG42;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG43;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG44;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG45;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG46;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG47;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG48;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG49;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG50;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG51;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG52;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG53;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG54;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG55;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG56;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG57;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG58;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG59;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG60;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG61;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG62;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG63;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG64;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG65;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG66;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG67;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG68;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG69;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG70;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG71;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG72;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG73;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG74;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG75;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG76;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG77;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG78;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG79;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG80;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG81;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG82;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG83;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG84;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG85;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG86;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG87;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG88;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG89;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG90;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG91;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG92;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG93;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG94;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG95;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG96;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG97;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG98;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG99;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOGSETN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRATOMICEGRESSBLOCKEDN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRCORN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRCPLABORTN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRCPLRDYN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRCPLTIMEOUTN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRCPLUNEXPECTN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRECRCN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRINTERNALCORN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRINTERNALUNCORN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRLOCKEDN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRMALFORMEDN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRMCBLOCKEDN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRNORECOVERYN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRPOISONEDN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRPOSTEDN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER32;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER33;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER34;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER35;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER36;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER37;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER38;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER39;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER40;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER41;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER42;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER43;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER44;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER45;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER46;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER47;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRURN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGFORCECOMMONCLOCKOFF;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGFORCEEXTENDEDSYNCON;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGFORCEMPS0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGFORCEMPS1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGFORCEMPS2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTASSERTN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTMMENABLE0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTMMENABLE1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTMMENABLE2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTMSIENABLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTMSIXENABLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTMSIXFM;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTRDYN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTSTATN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLASPMCONTROL0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLASPMCONTROL1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLAUTOBANDWIDTHINTEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLBANDWIDTHINTEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLCLOCKPMEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLCOMMONCLOCK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLEXTENDEDSYNC;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLHWAUTOWIDTHDIS;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLLINKDISABLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLRCB;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLRETRAINLINK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSAUTOBANDWIDTHSTATUS;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSBANDWIDTHSTATUS;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSCURRENTSPEED0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSCURRENTSPEED1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSDLLACTIVE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSLINKTRAINING;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSNEGOTIATEDWIDTH0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSNEGOTIATEDWIDTH1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSNEGOTIATEDWIDTH2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSNEGOTIATEDWIDTH3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTBYTEENN0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTBYTEENN1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTBYTEENN2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTBYTEENN3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTRDENN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTRDWRDONEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTWRENN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTWRREADONLYN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTWRRW1CASRWN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDASSERTINTA;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDASSERTINTB;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDASSERTINTC;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDASSERTINTD;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDDEASSERTINTA;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDDEASSERTINTB;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDDEASSERTINTC;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDDEASSERTINTD;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDERRCOR;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDERRFATAL;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDERRNONFATAL;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDPMASNAK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDPMETO;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDPMETOACK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDPMPME;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDSETSLOTPOWERLIMIT;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDUNLOCK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIECAPINTERRUPTMSGNUM0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIECAPINTERRUPTMSGNUM1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIECAPINTERRUPTMSGNUM2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIECAPINTERRUPTMSGNUM3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIECAPINTERRUPTMSGNUM4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIELINKSTATE0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIELINKSTATE1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIELINKSTATE2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMCSRPMEEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMCSRPMESTATUS;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMCSRPOWERSTATE0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMCSRPOWERSTATE1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMFORCESTATE0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMFORCESTATE1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMFORCESTATEENN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMHALTASPML0SN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMHALTASPML1N;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMRCVASREQL1N;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMRCVENTERL1N;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMRCVENTERL23N;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMRCVREQACKN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMSENDPMETON;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMTURNOFFOKN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMWAKEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGROOTCONTROLPMEINTEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGROOTCONTROLSYSERRCORRERREN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGROOTCONTROLSYSERRFATALERREN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGROOTCONTROLSYSERRNONFATALERREN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSLOTCONTROLELECTROMECHILCTLPULSE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTION;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONADDR0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONADDR1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONADDR2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONADDR3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONADDR4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONADDR5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONADDR6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONTYPE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRNPENDINGN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVCTCVCMAP0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVCTCVCMAP1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVCTCVCMAP2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVCTCVCMAP3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVCTCVCMAP4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVCTCVCMAP5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVCTCVCMAP6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CMRSTN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_CMSTICKYRSTN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGMODE0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGMODE1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRA;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRB;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRC;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRD;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRF;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRG;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRH;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRI;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRJ;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSUBMODE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA32;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA33;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA34;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA35;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA36;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA37;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA38;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA39;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA40;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA41;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA42;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA43;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA44;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA45;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA46;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA47;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA48;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA49;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA50;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA51;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA52;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA53;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA54;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA55;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA56;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA57;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA58;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA59;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA60;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA61;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA62;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA63;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB32;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB33;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB34;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB35;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB36;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB37;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB38;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB39;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB40;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB41;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB42;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB43;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB44;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB45;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB46;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB47;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB48;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB49;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB50;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB51;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB52;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB53;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB54;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB55;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB56;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB57;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB58;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB59;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB60;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB61;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB62;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB63;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DLRSTN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPCLK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPRDY;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_DRPWE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_FUNCLVLRSTN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2BADDLLPERR;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2BADTLPERR;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2LINKSTATUS0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2LINKSTATUS1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2LINKSTATUS2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2LINKSTATUS3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2LINKSTATUS4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2PROTOCOLERR;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2RECEIVERERR;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2REPLAYROERR;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2REPLAYTOERR;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2SENDASREQL1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2SENDENTERL1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2SENDENTERL23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2SENDPMACK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2SUSPENDNOW;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2SUSPENDOK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2TFCINIT1SEQ;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2TFCINIT2SEQ;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2TLPRCV;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LL2TXIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_LNKCLKEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA32;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA33;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA34;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA35;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA36;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA37;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA38;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA39;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA40;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA41;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA42;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA43;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA44;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA45;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA46;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA47;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA48;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA49;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA50;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA51;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA52;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA53;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA54;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA55;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA56;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA57;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA58;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA59;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA60;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA61;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA62;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA63;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA64;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA65;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA66;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA67;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXREN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA32;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA33;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA34;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA35;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA36;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA37;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA38;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA39;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA40;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA41;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA42;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA43;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA44;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA45;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA46;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA47;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA48;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA49;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA50;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA51;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA52;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA53;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA54;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA55;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA56;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA57;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA58;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA59;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA60;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA61;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA62;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA63;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA64;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA65;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA66;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA67;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA32;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA33;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA34;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA35;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA36;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA37;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA38;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA39;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA40;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA41;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA42;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA43;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA44;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA45;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA46;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA47;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA48;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA49;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA50;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA51;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA52;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA53;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA54;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA55;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA56;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA57;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA58;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA59;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA60;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA61;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA62;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA63;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA64;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA65;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA66;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA67;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA68;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXREN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA32;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA33;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA34;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA35;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA36;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA37;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA38;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA39;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA40;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA41;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA42;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA43;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA44;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA45;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA46;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA47;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA48;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA49;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA50;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA51;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA52;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA53;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA54;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA55;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA56;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA57;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA58;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA59;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA60;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA61;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA62;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA63;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA64;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA65;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA66;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA67;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA68;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPECLK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0CHANISALIGNED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0PHYSTATUS;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0POLARITY;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0STATUS0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0STATUS1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0STATUS2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0VALID;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1CHANISALIGNED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1PHYSTATUS;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1POLARITY;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1STATUS0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1STATUS1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1STATUS2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1VALID;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2CHANISALIGNED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2PHYSTATUS;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2POLARITY;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2STATUS0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2STATUS1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2STATUS2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2VALID;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3CHANISALIGNED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3PHYSTATUS;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3POLARITY;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3STATUS0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3STATUS1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3STATUS2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3VALID;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4CHANISALIGNED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4PHYSTATUS;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4POLARITY;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4STATUS0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4STATUS1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4STATUS2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4VALID;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5CHANISALIGNED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5PHYSTATUS;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5POLARITY;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5STATUS0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5STATUS1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5STATUS2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5VALID;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6CHANISALIGNED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6PHYSTATUS;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6POLARITY;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6STATUS0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6STATUS1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6STATUS2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6VALID;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7CHANISALIGNED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7PHYSTATUS;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7POLARITY;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7STATUS0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7STATUS1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7STATUS2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7VALID;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0COMPLIANCE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0POWERDOWN0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0POWERDOWN1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1COMPLIANCE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1POWERDOWN0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1POWERDOWN1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2COMPLIANCE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2POWERDOWN0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2POWERDOWN1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3COMPLIANCE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3POWERDOWN0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3POWERDOWN1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4COMPLIANCE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4POWERDOWN0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4POWERDOWN1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5COMPLIANCE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5POWERDOWN0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5POWERDOWN1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6COMPLIANCE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6POWERDOWN0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6POWERDOWN1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7CHARISK0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7CHARISK1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7COMPLIANCE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7ELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7POWERDOWN0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7POWERDOWN1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETXDEEMPH;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETXMARGIN0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETXMARGIN1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETXMARGIN2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETXRATE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETXRCVRDET;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETXRESET;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PL2DIRECTEDLSTATE0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PL2DIRECTEDLSTATE1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PL2DIRECTEDLSTATE2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PL2DIRECTEDLSTATE3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PL2DIRECTEDLSTATE4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PL2L0REQ;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PL2LINKUP;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PL2RECEIVERERR;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PL2RECOVERY;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PL2RXELECIDLE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PL2RXPMSTATE0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PL2RXPMSTATE1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PL2SUSPENDOK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGMODE0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGMODE1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGMODE2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDCHANGEDONE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLINKAUTON;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLINKCHANGE0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLINKCHANGE1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLINKSPEED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLINKWIDTH0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLINKWIDTH1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMNEW0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMNEW1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMNEW2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMNEW3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMNEW4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMNEW5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMNEWVLD;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMSTALL;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLDOWNSTREAMDEEMPHSOURCE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLINITIALLINKWIDTH0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLINITIALLINKWIDTH1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLINITIALLINKWIDTH2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLLANEREVERSALMODE0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLLANEREVERSALMODE1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLLINKGEN2CAP;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLLINKPARTNERGEN2SUPPORTED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLLINKUPCFGCAP;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLLTSSMSTATE0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLLTSSMSTATE1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLLTSSMSTATE2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLLTSSMSTATE3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLLTSSMSTATE4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLLTSSMSTATE5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLPHYLNKUPN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLRECEIVEDHOTRST;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLRSTN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLRXPMSTATE0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLRXPMSTATE1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLSELLNKRATE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLSELLNKWIDTH0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLSELLNKWIDTH1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLTRANSMITHOTRST;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLTXPMSTATE0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLTXPMSTATE1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLTXPMSTATE2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_PLUPSTREAMPREFERDEEMPH;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_RECEIVEDFUNCLVLRSTN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_SYSRSTN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ASPMSUSPENDCREDITCHECK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ASPMSUSPENDCREDITCHECKOK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ASPMSUSPENDREQ;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRFCPE;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR32;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR33;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR34;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR35;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR36;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR37;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR38;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR39;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR40;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR41;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR42;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR43;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR44;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR45;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR46;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR47;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR48;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR49;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR50;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR51;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR52;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR53;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR54;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR55;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR56;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR57;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR58;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR59;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR60;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR61;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR62;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR63;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRMALFORMED;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRRXOVERFLOW;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2PPMSUSPENDOK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TL2PPMSUSPENDREQ;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TLRSTN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCSEL0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCSEL1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCSEL2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNLNKUP;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD100;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD101;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD102;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD103;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD104;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD105;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD106;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD107;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD108;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD109;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD110;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD111;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD112;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD113;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD114;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD115;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD116;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD117;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD118;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD119;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD120;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD121;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD122;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD123;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD124;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD125;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD126;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD127;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD32;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD33;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD34;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD35;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD36;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD37;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD38;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD39;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD40;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD41;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD42;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD43;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD44;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD45;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD46;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD47;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD48;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD49;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD50;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD51;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD52;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD53;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD54;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD55;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD56;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD57;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD58;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD59;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD60;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD61;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD62;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD63;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD64;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD65;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD66;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD67;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD68;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD69;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD70;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD71;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD72;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD73;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD74;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD75;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD76;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD77;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD78;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD79;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD80;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD81;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD82;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD83;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD84;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD85;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD86;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD87;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD88;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD89;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD90;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD91;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD92;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD93;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD94;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD95;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD96;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD97;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD98;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD99;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA32;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA33;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA34;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA35;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA36;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA37;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA38;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA39;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA40;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA41;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA42;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA43;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA44;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA45;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA46;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA47;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA48;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA49;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA50;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA51;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA52;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA53;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA54;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA55;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA56;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA57;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA58;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA59;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA60;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA61;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA62;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA63;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPSRCRDY0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPSRCRDY1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDSTRDY;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRECRCERR;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNREOF;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRERRFWD;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRFCPRET;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRNPOK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRNPREQ;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRREM0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRREM1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRSOF;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRSRCDSC;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRSRCRDY;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTBUFAV0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTBUFAV1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTBUFAV2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTBUFAV3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTBUFAV4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTBUFAV5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTCFGGNT;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTCFGREQ;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD100;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD101;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD102;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD103;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD104;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD105;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD106;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD107;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD108;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD109;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD110;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD111;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD112;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD113;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD114;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD115;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD116;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD117;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD118;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD119;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD120;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD121;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD122;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD123;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD124;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD125;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD126;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD127;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD32;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD33;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD34;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD35;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD36;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD37;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD38;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD39;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD40;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD41;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD42;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD43;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD44;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD45;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD46;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD47;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD48;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD49;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD50;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD51;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD52;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD53;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD54;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD55;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD56;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD57;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD58;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD59;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD60;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD61;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD62;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD63;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD64;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD65;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD66;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD67;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD68;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD69;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD70;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD71;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD72;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD73;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD74;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD75;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD76;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD77;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD78;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD79;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD80;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD81;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD82;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD83;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD84;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD85;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD86;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD87;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD88;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD89;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD90;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD91;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD92;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD93;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD94;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD95;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD96;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD97;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD98;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD99;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA10;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA11;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA12;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA13;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA14;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA15;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA16;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA17;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA18;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA19;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA20;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA21;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA22;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA23;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA24;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA25;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA26;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA27;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA28;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA29;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA30;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA31;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA4;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA5;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA6;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA7;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA8;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA9;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDSTRDY;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPSRCRDY;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDSTRDY0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDSTRDY1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDSTRDY2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDSTRDY3;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTECRCGEN;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTEOF;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTERRDROP;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTERRFWD;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTREM0;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTREM1;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTSOF;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTSRCDSC;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTSRCRDY;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTSTR;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_USERCLK;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_USERCLK2;
  wire [0:0] PCIE_BOT_X71Y115_PCIE_X0Y0_USERRSTN;
  wire [0:0] RIOB33_X43Y31_IOB_X1Y32_O;
  wire [0:0] RIOB33_X43Y37_IOB_X1Y37_O;
  wire [0:0] RIOB33_X43Y37_IOB_X1Y38_O;
  wire [0:0] RIOB33_X43Y39_IOB_X1Y39_I;
  wire [0:0] RIOB33_X43Y39_IOB_X1Y40_I;
  wire [0:0] RIOB33_X43Y43_IOB_X1Y43_I;
  wire [0:0] RIOB33_X43Y43_IOB_X1Y44_I;
  wire [0:0] RIOB33_X43Y45_IOB_X1Y45_I;
  wire [0:0] RIOB33_X43Y45_IOB_X1Y46_I;
  wire [0:0] RIOB33_X43Y47_IOB_X1Y47_I;
  wire [0:0] RIOB33_X43Y47_IOB_X1Y48_I;
  wire [0:0] RIOB33_X43Y61_IOB_X1Y61_O;
  wire [0:0] RIOB33_X43Y75_IOB_X1Y75_O;
  wire [0:0] RIOB33_X43Y75_IOB_X1Y76_O;
  wire [0:0] RIOB33_X43Y87_IOB_X1Y87_O;
  wire [0:0] RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_D1;
  wire [0:0] RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_OQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_T1;
  wire [0:0] RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_TQ;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_D;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_O;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_D;
  wire [0:0] RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_O;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_D1;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_OQ;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_T1;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_TQ;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_D1;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_OQ;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_T1;
  wire [0:0] RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_TQ;
  wire [0:0] RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_D1;
  wire [0:0] RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_OQ;
  wire [0:0] RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_T1;
  wire [0:0] RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_TQ;
  wire [0:0] RIOI3_X43Y39_ILOGIC_X1Y39_D;
  wire [0:0] RIOI3_X43Y39_ILOGIC_X1Y39_O;
  wire [0:0] RIOI3_X43Y39_ILOGIC_X1Y40_D;
  wire [0:0] RIOI3_X43Y39_ILOGIC_X1Y40_O;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y45_D;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y45_O;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y46_D;
  wire [0:0] RIOI3_X43Y45_ILOGIC_X1Y46_O;
  wire [0:0] RIOI3_X43Y47_ILOGIC_X1Y47_D;
  wire [0:0] RIOI3_X43Y47_ILOGIC_X1Y47_O;
  wire [0:0] RIOI3_X43Y47_ILOGIC_X1Y48_D;
  wire [0:0] RIOI3_X43Y47_ILOGIC_X1Y48_O;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_D1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_OQ;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_T1;
  wire [0:0] RIOI3_X43Y61_OLOGIC_X1Y61_TQ;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y75_D1;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y75_OQ;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y75_T1;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y75_TQ;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y76_D1;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y76_OQ;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y76_T1;
  wire [0:0] RIOI3_X43Y75_OLOGIC_X1Y76_TQ;


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y1_OBUF (
.I(LIOB33_X0Y5_IOB_X0Y6_I),
.O(led[7])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y1_IOB_X0Y2_OBUF (
.I(RIOB33_X43Y39_IOB_X1Y40_I),
.O(led[8])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y3_IOB_X0Y3_OBUF (
.I(PCIE_BOT_X71Y115_PCIE_X0Y0_DRPRDY),
.O(led[0])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y3_IOB_X0Y4_OBUF (
.I(LIOB33_X0Y7_IOB_X0Y8_I),
.O(led[5])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y5_IOB_X0Y5_IBUF (
.I(sw[6]),
.O(LIOB33_X0Y5_IOB_X0Y5_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y5_IOB_X0Y6_IBUF (
.I(sw[7]),
.O(LIOB33_X0Y5_IOB_X0Y6_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y7_IOB_X0Y7_IBUF (
.I(sw[4]),
.O(LIOB33_X0Y7_IOB_X0Y7_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y7_IOB_X0Y8_IBUF (
.I(sw[5]),
.O(LIOB33_X0Y7_IOB_X0Y8_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y9_IOB_X0Y9_IBUF (
.I(sw[3]),
.O(LIOB33_X0Y9_IOB_X0Y9_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y9_IOB_X0Y10_IBUF (
.I(sw[2]),
.O(LIOB33_X0Y9_IOB_X0Y10_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y11_IOB_X0Y11_IBUF (
.I(sw[0]),
.O(LIOB33_X0Y11_IOB_X0Y11_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y11_IOB_X0Y12_IBUF (
.I(sw[1]),
.O(LIOB33_X0Y11_IOB_X0Y12_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y17_IOB_X0Y18_OBUF (
.I(LIOB33_X0Y7_IOB_X0Y7_I),
.O(led[4])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y19_IOB_X0Y19_OBUF (
.I(LIOB33_X0Y9_IOB_X0Y9_I),
.O(led[3])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y19_IOB_X0Y20_OBUF (
.I(LIOB33_X0Y9_IOB_X0Y10_I),
.O(led[2])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y43_IOB_X0Y43_OBUF (
.I(LIOB33_X0Y11_IOB_X0Y12_I),
.O(led[1])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y111_IOB_X0Y111_OBUF (
.I(LIOB33_X0Y111_IOB_X0Y112_I),
.O(tx)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y111_IOB_X0Y112_IBUF (
.I(rx),
.O(LIOB33_X0Y111_IOB_X0Y112_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_SING_X0Y0_IOB_X0Y0_OBUF (
.I(LIOB33_X0Y5_IOB_X0Y5_I),
.O(led[6])
  );


  (* KEEP, DONT_TOUCH, BEL = "PCIE_2_1" *)
  PCIE_2_1 #(
    .AER_BASE_PTR(12'b000000000000),
    .AER_CAP_ECRC_CHECK_CAPABLE("FALSE"),
    .AER_CAP_ECRC_GEN_CAPABLE("FALSE"),
    .AER_CAP_ID(16'b0000000000000000),
    .AER_CAP_MULTIHEADER("FALSE"),
    .AER_CAP_NEXTPTR(12'b000000000000),
    .AER_CAP_ON("FALSE"),
    .AER_CAP_OPTIONAL_ERR_SUPPORT(24'b000000000000000000000000),
    .AER_CAP_PERMIT_ROOTERR_UPDATE("FALSE"),
    .AER_CAP_VERSION(4'b0000),
    .ALLOW_X8_GEN2("FALSE"),
    .BAR0(32'b00000000000000000000000000000000),
    .BAR1(32'b00000000000000000000000000000000),
    .BAR2(32'b00000000000000000000000000000000),
    .BAR3(32'b00000000000000000000000000000000),
    .BAR4(32'b00000000000000000000000000000000),
    .BAR5(32'b00000000000000000000000000000000),
    .CAPABILITIES_PTR(8'b00000000),
    .CARDBUS_CIS_POINTER(32'b00000000000000000000000000000000),
    .CFG_ECRC_ERR_CPLSTAT(2'b00),
    .CLASS_CODE(24'b000000000000000000000000),
    .CMD_INTX_IMPLEMENTED("FALSE"),
    .CPL_TIMEOUT_DISABLE_SUPPORTED("FALSE"),
    .CPL_TIMEOUT_RANGES_SUPPORTED(4'b0000),
    .CRM_MODULE_RSTS(7'b0000000),
    .DEV_CAP2_ARI_FORWARDING_SUPPORTED("FALSE"),
    .DEV_CAP2_ATOMICOP32_COMPLETER_SUPPORTED("FALSE"),
    .DEV_CAP2_ATOMICOP64_COMPLETER_SUPPORTED("FALSE"),
    .DEV_CAP2_ATOMICOP_ROUTING_SUPPORTED("FALSE"),
    .DEV_CAP2_CAS128_COMPLETER_SUPPORTED("FALSE"),
    .DEV_CAP2_ENDEND_TLP_PREFIX_SUPPORTED("FALSE"),
    .DEV_CAP2_EXTENDED_FMT_FIELD_SUPPORTED("FALSE"),
    .DEV_CAP2_LTR_MECHANISM_SUPPORTED("FALSE"),
    .DEV_CAP2_MAX_ENDEND_TLP_PREFIXES(2'b00),
    .DEV_CAP2_NO_RO_ENABLED_PRPR_PASSING("FALSE"),
    .DEV_CAP2_TPH_COMPLETER_SUPPORTED(2'b00),
    .DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE("FALSE"),
    .DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE("FALSE"),
    .DEV_CAP_ENDPOINT_L0S_LATENCY(3'b000),
    .DEV_CAP_ENDPOINT_L1_LATENCY(3'b000),
    .DEV_CAP_EXT_TAG_SUPPORTED("FALSE"),
    .DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE("FALSE"),
    .DEV_CAP_MAX_PAYLOAD_SUPPORTED(3'b000),
    .DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT(2'b00),
    .DEV_CAP_ROLE_BASED_ERROR("FALSE"),
    .DEV_CAP_RSVD_14_12(3'b000),
    .DEV_CAP_RSVD_17_16(2'b00),
    .DEV_CAP_RSVD_31_29(3'b000),
    .DEV_CONTROL_AUX_POWER_SUPPORTED("FALSE"),
    .DEV_CONTROL_EXT_TAG_DEFAULT("FALSE"),
    .DISABLE_ASPM_L1_TIMER("FALSE"),
    .DISABLE_BAR_FILTERING("FALSE"),
    .DISABLE_ERR_MSG("FALSE"),
    .DISABLE_ID_CHECK("FALSE"),
    .DISABLE_LANE_REVERSAL("FALSE"),
    .DISABLE_LOCKED_FILTER("FALSE"),
    .DISABLE_PPM_FILTER("FALSE"),
    .DISABLE_RX_POISONED_RESP("FALSE"),
    .DISABLE_RX_TC_FILTER("FALSE"),
    .DISABLE_SCRAMBLING("FALSE"),
    .DNSTREAM_LINK_NUM(8'b00000000),
    .DSN_BASE_PTR(12'b000000000000),
    .DSN_CAP_ID(16'b0000000000000000),
    .DSN_CAP_NEXTPTR(12'b000000000000),
    .DSN_CAP_ON("FALSE"),
    .DSN_CAP_VERSION(4'b0000),
    .ENABLE_MSG_ROUTE(11'b00000000000),
    .ENABLE_RX_TD_ECRC_TRIM("FALSE"),
    .ENDEND_TLP_PREFIX_FORWARDING_SUPPORTED("FALSE"),
    .ENTER_RVRY_EI_L0("FALSE"),
    .EXIT_LOOPBACK_ON_EI("FALSE"),
    .EXPANSION_ROM(32'b00000000000000000000000000000000),
    .EXT_CFG_CAP_PTR(6'b000000),
    .EXT_CFG_XP_CAP_PTR(10'b0000000000),
    .HEADER_TYPE(8'b00000000),
    .INFER_EI(5'b00000),
    .INTERRUPT_PIN(8'b00000000),
    .INTERRUPT_STAT_AUTO("FALSE"),
    .IS_SWITCH("FALSE"),
    .LAST_CONFIG_DWORD(10'b0000000000),
    .LINK_CAP_ASPM_OPTIONALITY("FALSE"),
    .LINK_CAP_ASPM_SUPPORT(2'b00),
    .LINK_CAP_CLOCK_POWER_MANAGEMENT("FALSE"),
    .LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP("FALSE"),
    .LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1(3'b000),
    .LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2(3'b000),
    .LINK_CAP_L0S_EXIT_LATENCY_GEN1(3'b000),
    .LINK_CAP_L0S_EXIT_LATENCY_GEN2(3'b000),
    .LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1(3'b000),
    .LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2(3'b000),
    .LINK_CAP_L1_EXIT_LATENCY_GEN1(3'b000),
    .LINK_CAP_L1_EXIT_LATENCY_GEN2(3'b000),
    .LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP("FALSE"),
    .LINK_CAP_MAX_LINK_SPEED(4'b0000),
    .LINK_CAP_MAX_LINK_WIDTH(6'b001000),
    .LINK_CAP_RSVD_23(1'b0),
    .LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE("FALSE"),
    .LINK_CONTROL_RCB(1'b0),
    .LINK_CTRL2_DEEMPHASIS("FALSE"),
    .LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE("FALSE"),
    .LINK_CTRL2_TARGET_LINK_SPEED(4'b0000),
    .LINK_STATUS_SLOT_CLOCK_CONFIG("FALSE"),
    .LL_ACK_TIMEOUT(15'b000000000000000),
    .LL_ACK_TIMEOUT_EN("FALSE"),
    .LL_ACK_TIMEOUT_FUNC(2'b00),
    .LL_REPLAY_TIMEOUT(15'b000000000000000),
    .LL_REPLAY_TIMEOUT_EN("FALSE"),
    .LL_REPLAY_TIMEOUT_FUNC(2'b00),
    .LTSSM_MAX_LINK_WIDTH(6'b000000),
    .MPS_FORCE("FALSE"),
    .MSIX_BASE_PTR(8'b00000000),
    .MSIX_CAP_ID(8'b00000000),
    .MSIX_CAP_NEXTPTR(8'b00000000),
    .MSIX_CAP_ON("FALSE"),
    .MSIX_CAP_PBA_BIR(3'b000),
    .MSIX_CAP_PBA_OFFSET(29'b00000000000000000000000000000),
    .MSIX_CAP_TABLE_BIR(3'b000),
    .MSIX_CAP_TABLE_OFFSET(29'b00000000000000000000000000000),
    .MSIX_CAP_TABLE_SIZE(11'b00000000000),
    .MSI_BASE_PTR(8'b00000000),
    .MSI_CAP_64_BIT_ADDR_CAPABLE("FALSE"),
    .MSI_CAP_ID(8'b00000000),
    .MSI_CAP_MULTIMSGCAP(3'b000),
    .MSI_CAP_MULTIMSG_EXTENSION(1'b0),
    .MSI_CAP_NEXTPTR(8'b00000000),
    .MSI_CAP_ON("FALSE"),
    .MSI_CAP_PER_VECTOR_MASKING_CAPABLE("FALSE"),
    .N_FTS_COMCLK_GEN1(8'b11111111),
    .N_FTS_COMCLK_GEN2(8'b11111111),
    .N_FTS_GEN1(8'b11111111),
    .N_FTS_GEN2(8'b11111111),
    .PCIE_BASE_PTR(8'b00000000),
    .PCIE_CAP_CAPABILITY_ID(8'b00000000),
    .PCIE_CAP_CAPABILITY_VERSION(4'b0000),
    .PCIE_CAP_DEVICE_PORT_TYPE(4'b0000),
    .PCIE_CAP_NEXTPTR(8'b00000000),
    .PCIE_CAP_ON("FALSE"),
    .PCIE_CAP_RSVD_15_14(2'b00),
    .PCIE_CAP_SLOT_IMPLEMENTED("FALSE"),
    .PCIE_REVISION(4'b0010),
    .PL_AUTO_CONFIG(3'b000),
    .PL_FAST_TRAIN("FALSE"),
    .PM_ASPML0S_TIMEOUT(15'b000000000000000),
    .PM_ASPML0S_TIMEOUT_EN("FALSE"),
    .PM_ASPML0S_TIMEOUT_FUNC(2'b00),
    .PM_ASPM_FASTEXIT("FALSE"),
    .PM_BASE_PTR(8'b00000000),
    .PM_CAP_AUXCURRENT(3'b000),
    .PM_CAP_D1SUPPORT("FALSE"),
    .PM_CAP_D2SUPPORT("FALSE"),
    .PM_CAP_DSI("FALSE"),
    .PM_CAP_ID(8'b00000000),
    .PM_CAP_NEXTPTR(8'b00000000),
    .PM_CAP_ON("FALSE"),
    .PM_CAP_PMESUPPORT(5'b00000),
    .PM_CAP_PME_CLOCK("FALSE"),
    .PM_CAP_RSVD_04(1'b0),
    .PM_CAP_VERSION(3'b011),
    .PM_CSR_B2B3("FALSE"),
    .PM_CSR_BPCCEN("FALSE"),
    .PM_CSR_NOSOFTRST("FALSE"),
    .PM_DATA0(8'b00000000),
    .PM_DATA1(8'b00000000),
    .PM_DATA2(8'b00000000),
    .PM_DATA3(8'b00000000),
    .PM_DATA4(8'b00000000),
    .PM_DATA5(8'b00000000),
    .PM_DATA6(8'b00000000),
    .PM_DATA7(8'b00000000),
    .PM_DATA_SCALE0(2'b00),
    .PM_DATA_SCALE1(2'b00),
    .PM_DATA_SCALE2(2'b00),
    .PM_DATA_SCALE3(2'b00),
    .PM_DATA_SCALE4(2'b00),
    .PM_DATA_SCALE5(2'b00),
    .PM_DATA_SCALE6(2'b00),
    .PM_DATA_SCALE7(2'b00),
    .PM_MF("FALSE"),
    .RBAR_BASE_PTR(12'b000000000000),
    .RBAR_CAP_CONTROL_ENCODEDBAR0(5'b00000),
    .RBAR_CAP_CONTROL_ENCODEDBAR1(5'b00000),
    .RBAR_CAP_CONTROL_ENCODEDBAR2(5'b00000),
    .RBAR_CAP_CONTROL_ENCODEDBAR3(5'b00000),
    .RBAR_CAP_CONTROL_ENCODEDBAR4(5'b00000),
    .RBAR_CAP_CONTROL_ENCODEDBAR5(5'b00000),
    .RBAR_CAP_ID(16'b0000000000000000),
    .RBAR_CAP_INDEX0(3'b000),
    .RBAR_CAP_INDEX1(3'b000),
    .RBAR_CAP_INDEX2(3'b000),
    .RBAR_CAP_INDEX3(3'b000),
    .RBAR_CAP_INDEX4(3'b000),
    .RBAR_CAP_INDEX5(3'b000),
    .RBAR_CAP_NEXTPTR(12'b000000000000),
    .RBAR_CAP_ON("FALSE"),
    .RBAR_CAP_SUP0(32'b00000000000000000000000000000000),
    .RBAR_CAP_SUP1(32'b00000000000000000000000000000000),
    .RBAR_CAP_SUP2(32'b00000000000000000000000000000000),
    .RBAR_CAP_SUP3(32'b00000000000000000000000000000000),
    .RBAR_CAP_SUP4(32'b00000000000000000000000000000000),
    .RBAR_CAP_SUP5(32'b00000000000000000000000000000000),
    .RBAR_CAP_VERSION(4'b0000),
    .RBAR_NUM(3'b000),
    .RECRC_CHK(2'b00),
    .RECRC_CHK_TRIM("FALSE"),
    .ROOT_CAP_CRS_SW_VISIBILITY("FALSE"),
    .RP_AUTO_SPD(2'b00),
    .RP_AUTO_SPD_LOOPCNT(5'b00000),
    .SELECT_DLL_IF("FALSE"),
    .SLOT_CAP_ATT_BUTTON_PRESENT("FALSE"),
    .SLOT_CAP_ATT_INDICATOR_PRESENT("FALSE"),
    .SLOT_CAP_ELEC_INTERLOCK_PRESENT("FALSE"),
    .SLOT_CAP_HOTPLUG_CAPABLE("FALSE"),
    .SLOT_CAP_HOTPLUG_SURPRISE("FALSE"),
    .SLOT_CAP_MRL_SENSOR_PRESENT("FALSE"),
    .SLOT_CAP_NO_CMD_COMPLETED_SUPPORT("FALSE"),
    .SLOT_CAP_PHYSICAL_SLOT_NUM(13'b0000000000000),
    .SLOT_CAP_POWER_CONTROLLER_PRESENT("FALSE"),
    .SLOT_CAP_POWER_INDICATOR_PRESENT("FALSE"),
    .SLOT_CAP_SLOT_POWER_LIMIT_SCALE(2'b00),
    .SLOT_CAP_SLOT_POWER_LIMIT_VALUE(8'b00000000),
    .SPARE_BIT0(1'b0),
    .SPARE_BIT1(1'b0),
    .SPARE_BIT2(1'b0),
    .SPARE_BIT3(1'b0),
    .SPARE_BIT4(1'b0),
    .SPARE_BIT5(1'b0),
    .SPARE_BIT6(1'b0),
    .SPARE_BIT7(1'b0),
    .SPARE_BIT8(1'b0),
    .SPARE_BYTE0(8'b00000000),
    .SPARE_BYTE1(8'b00000000),
    .SPARE_BYTE2(8'b00000000),
    .SPARE_BYTE3(8'b00000000),
    .SPARE_WORD0(32'b00000000000000000000000000000000),
    .SPARE_WORD1(32'b00000000000000000000000000000000),
    .SPARE_WORD2(32'b00000000000000000000000000000000),
    .SPARE_WORD3(32'b00000000000000000000000000000000),
    .SSL_MESSAGE_AUTO("FALSE"),
    .TECRC_EP_INV("FALSE"),
    .TL_RBYPASS("FALSE"),
    .TL_RX_RAM_RADDR_LATENCY(1'b0),
    .TL_RX_RAM_RDATA_LATENCY(2'b01),
    .TL_RX_RAM_WRITE_LATENCY(1'b0),
    .TL_TFC_DISABLE("FALSE"),
    .TL_TX_CHECKS_DISABLE("FALSE"),
    .TL_TX_RAM_RADDR_LATENCY(1'b0),
    .TL_TX_RAM_RDATA_LATENCY(2'b01),
    .TL_TX_RAM_WRITE_LATENCY(1'b0),
    .TRN_DW("FALSE"),
    .TRN_NP_FC("FALSE"),
    .UPCONFIG_CAPABLE("FALSE"),
    .UPSTREAM_FACING("FALSE"),
    .UR_ATOMIC("FALSE"),
    .UR_CFG1("FALSE"),
    .UR_INV_REQ("FALSE"),
    .UR_PRS_RESPONSE("FALSE"),
    .USER_CLK2_DIV2("FALSE"),
    .USER_CLK_FREQ(3'b000),
    .USE_RID_PINS("FALSE"),
    .VC0_CPL_INFINITE("FALSE"),
    .VC0_RX_RAM_LIMIT(13'b0000000000000),
    .VC0_TOTAL_CREDITS_CD(11'b00000000000),
    .VC0_TOTAL_CREDITS_CH(7'b0100100),
    .VC0_TOTAL_CREDITS_NPD(11'b00000000000),
    .VC0_TOTAL_CREDITS_NPH(7'b0001100),
    .VC0_TOTAL_CREDITS_PD(11'b00000000000),
    .VC0_TOTAL_CREDITS_PH(7'b0100000),
    .VC0_TX_LASTPACKET(5'b00000),
    .VC_BASE_PTR(12'b000000000000),
    .VC_CAP_ID(16'b0000000000000000),
    .VC_CAP_NEXTPTR(12'b000000000000),
    .VC_CAP_ON("FALSE"),
    .VC_CAP_REJECT_SNOOP_TRANSACTIONS("FALSE"),
    .VC_CAP_VERSION(4'b0000),
    .VSEC_BASE_PTR(12'b000000000000),
    .VSEC_CAP_HDR_ID(16'b0000000000000000),
    .VSEC_CAP_HDR_LENGTH(12'b000000000000),
    .VSEC_CAP_HDR_REVISION(4'b0000),
    .VSEC_CAP_ID(16'b0000000000000000),
    .VSEC_CAP_IS_LINK_VISIBLE("FALSE"),
    .VSEC_CAP_NEXTPTR(12'b000000000000),
    .VSEC_CAP_ON("FALSE"),
    .VSEC_CAP_VERSION(4'b0000)
  ) PCIE_BOT_X71Y115_PCIE_X0Y0_PCIE_2_1 (
.CFGAERECRCCHECKEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERECRCCHECKEN),
.CFGAERECRCGENEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERECRCGENEN),
.CFGAERINTERRUPTMSGNUM({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CFGAERROOTERRCORRERRRECEIVED(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERROOTERRCORRERRRECEIVED),
.CFGAERROOTERRCORRERRREPORTINGEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERROOTERRCORRERRREPORTINGEN),
.CFGAERROOTERRFATALERRRECEIVED(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERROOTERRFATALERRRECEIVED),
.CFGAERROOTERRFATALERRREPORTINGEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERROOTERRFATALERRREPORTINGEN),
.CFGAERROOTERRNONFATALERRRECEIVED(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERROOTERRNONFATALERRRECEIVED),
.CFGAERROOTERRNONFATALERRREPORTINGEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERROOTERRNONFATALERRREPORTINGEN),
.CFGBRIDGESERREN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGBRIDGESERREN),
.CFGCOMMANDBUSMASTERENABLE(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGCOMMANDBUSMASTERENABLE),
.CFGCOMMANDINTERRUPTDISABLE(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGCOMMANDINTERRUPTDISABLE),
.CFGCOMMANDIOENABLE(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGCOMMANDIOENABLE),
.CFGCOMMANDMEMENABLE(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGCOMMANDMEMENABLE),
.CFGCOMMANDSERREN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGCOMMANDSERREN),
.CFGDEVCONTROL2ARIFORWARDEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2ARIFORWARDEN),
.CFGDEVCONTROL2ATOMICEGRESSBLOCK(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2ATOMICEGRESSBLOCK),
.CFGDEVCONTROL2ATOMICREQUESTEREN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2ATOMICREQUESTEREN),
.CFGDEVCONTROL2CPLTIMEOUTDIS(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2CPLTIMEOUTDIS),
.CFGDEVCONTROL2CPLTIMEOUTVAL({PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2CPLTIMEOUTVAL3, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2CPLTIMEOUTVAL2, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2CPLTIMEOUTVAL1, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2CPLTIMEOUTVAL0}),
.CFGDEVCONTROL2IDOCPLEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2IDOCPLEN),
.CFGDEVCONTROL2IDOREQEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2IDOREQEN),
.CFGDEVCONTROL2LTREN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2LTREN),
.CFGDEVCONTROL2TLPPREFIXBLOCK(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROL2TLPPREFIXBLOCK),
.CFGDEVCONTROLAUXPOWEREN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLAUXPOWEREN),
.CFGDEVCONTROLCORRERRREPORTINGEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLCORRERRREPORTINGEN),
.CFGDEVCONTROLENABLERO(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLENABLERO),
.CFGDEVCONTROLEXTTAGEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLEXTTAGEN),
.CFGDEVCONTROLFATALERRREPORTINGEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLFATALERRREPORTINGEN),
.CFGDEVCONTROLMAXPAYLOAD({PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLMAXPAYLOAD2, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLMAXPAYLOAD1, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLMAXPAYLOAD0}),
.CFGDEVCONTROLMAXREADREQ({PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLMAXREADREQ2, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLMAXREADREQ1, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLMAXREADREQ0}),
.CFGDEVCONTROLNONFATALREPORTINGEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLNONFATALREPORTINGEN),
.CFGDEVCONTROLNOSNOOPEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLNOSNOOPEN),
.CFGDEVCONTROLPHANTOMEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLPHANTOMEN),
.CFGDEVCONTROLURERRREPORTINGEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVCONTROLURERRREPORTINGEN),
.CFGDEVID({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CFGDEVSTATUSCORRERRDETECTED(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVSTATUSCORRERRDETECTED),
.CFGDEVSTATUSFATALERRDETECTED(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVSTATUSFATALERRDETECTED),
.CFGDEVSTATUSNONFATALERRDETECTED(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVSTATUSNONFATALERRDETECTED),
.CFGDEVSTATUSURDETECTED(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVSTATUSURDETECTED),
.CFGDSBUSNUMBER({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CFGDSDEVICENUMBER({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CFGDSFUNCTIONNUMBER({1'b0, 1'b0, 1'b0}),
.CFGDSN({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CFGERRACSN(1'b0),
.CFGERRAERHEADERLOG({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CFGERRAERHEADERLOGSETN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOGSETN),
.CFGERRATOMICEGRESSBLOCKEDN(1'b0),
.CFGERRCORN(1'b0),
.CFGERRCPLABORTN(1'b0),
.CFGERRCPLRDYN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRCPLRDYN),
.CFGERRCPLTIMEOUTN(1'b0),
.CFGERRCPLUNEXPECTN(1'b0),
.CFGERRECRCN(1'b0),
.CFGERRINTERNALCORN(1'b0),
.CFGERRINTERNALUNCORN(1'b0),
.CFGERRLOCKEDN(1'b0),
.CFGERRMALFORMEDN(1'b0),
.CFGERRMCBLOCKEDN(1'b0),
.CFGERRNORECOVERYN(1'b0),
.CFGERRPOISONEDN(1'b0),
.CFGERRPOSTEDN(1'b0),
.CFGERRTLPCPLHEADER({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CFGERRURN(1'b0),
.CFGFORCECOMMONCLOCKOFF(1'b0),
.CFGFORCEEXTENDEDSYNCON(1'b0),
.CFGFORCEMPS({1'b0, 1'b0, 1'b0}),
.CFGINTERRUPTASSERTN(1'b0),
.CFGINTERRUPTDI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CFGINTERRUPTDO({PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO7, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO6, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO5, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO4, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO3, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO2, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO1, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDO0}),
.CFGINTERRUPTMMENABLE({PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTMMENABLE2, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTMMENABLE1, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTMMENABLE0}),
.CFGINTERRUPTMSIENABLE(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTMSIENABLE),
.CFGINTERRUPTMSIXENABLE(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTMSIXENABLE),
.CFGINTERRUPTMSIXFM(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTMSIXFM),
.CFGINTERRUPTN(1'b0),
.CFGINTERRUPTRDYN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTRDYN),
.CFGINTERRUPTSTATN(1'b0),
.CFGLINKCONTROLASPMCONTROL({PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLASPMCONTROL1, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLASPMCONTROL0}),
.CFGLINKCONTROLAUTOBANDWIDTHINTEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLAUTOBANDWIDTHINTEN),
.CFGLINKCONTROLBANDWIDTHINTEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLBANDWIDTHINTEN),
.CFGLINKCONTROLCLOCKPMEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLCLOCKPMEN),
.CFGLINKCONTROLCOMMONCLOCK(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLCOMMONCLOCK),
.CFGLINKCONTROLEXTENDEDSYNC(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLEXTENDEDSYNC),
.CFGLINKCONTROLHWAUTOWIDTHDIS(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLHWAUTOWIDTHDIS),
.CFGLINKCONTROLLINKDISABLE(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLLINKDISABLE),
.CFGLINKCONTROLRCB(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLRCB),
.CFGLINKCONTROLRETRAINLINK(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKCONTROLRETRAINLINK),
.CFGLINKSTATUSAUTOBANDWIDTHSTATUS(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSAUTOBANDWIDTHSTATUS),
.CFGLINKSTATUSBANDWIDTHSTATUS(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSBANDWIDTHSTATUS),
.CFGLINKSTATUSCURRENTSPEED({PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSCURRENTSPEED1, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSCURRENTSPEED0}),
.CFGLINKSTATUSDLLACTIVE(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSDLLACTIVE),
.CFGLINKSTATUSLINKTRAINING(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSLINKTRAINING),
.CFGLINKSTATUSNEGOTIATEDWIDTH({PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSNEGOTIATEDWIDTH3, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSNEGOTIATEDWIDTH2, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSNEGOTIATEDWIDTH1, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGLINKSTATUSNEGOTIATEDWIDTH0}),
.CFGMGMTBYTEENN({1'b0, 1'b0, 1'b0, 1'b0}),
.CFGMGMTDI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CFGMGMTDO({PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO31, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO30, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO29, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO28, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO27, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO26, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO25, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO24, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO23, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO22, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO21, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO20, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO19, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO18, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO17, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO16, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO15, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO14, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO13, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO12, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO11, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO10, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO9, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO8, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO7, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO6, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO5, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO4, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO3, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO2, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO1, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDO0}),
.CFGMGMTDWADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CFGMGMTRDENN(1'b0),
.CFGMGMTRDWRDONEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTRDWRDONEN),
.CFGMGMTWRENN(1'b0),
.CFGMGMTWRREADONLYN(1'b0),
.CFGMGMTWRRW1CASRWN(1'b0),
.CFGMSGDATA({PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA15, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA14, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA13, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA12, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA11, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA10, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA9, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA8, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA7, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA6, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA5, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA4, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA3, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA2, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA1, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGDATA0}),
.CFGMSGRECEIVED(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVED),
.CFGMSGRECEIVEDASSERTINTA(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDASSERTINTA),
.CFGMSGRECEIVEDASSERTINTB(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDASSERTINTB),
.CFGMSGRECEIVEDASSERTINTC(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDASSERTINTC),
.CFGMSGRECEIVEDASSERTINTD(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDASSERTINTD),
.CFGMSGRECEIVEDDEASSERTINTA(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDDEASSERTINTA),
.CFGMSGRECEIVEDDEASSERTINTB(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDDEASSERTINTB),
.CFGMSGRECEIVEDDEASSERTINTC(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDDEASSERTINTC),
.CFGMSGRECEIVEDDEASSERTINTD(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDDEASSERTINTD),
.CFGMSGRECEIVEDERRCOR(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDERRCOR),
.CFGMSGRECEIVEDERRFATAL(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDERRFATAL),
.CFGMSGRECEIVEDERRNONFATAL(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDERRNONFATAL),
.CFGMSGRECEIVEDPMASNAK(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDPMASNAK),
.CFGMSGRECEIVEDPMETO(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDPMETO),
.CFGMSGRECEIVEDPMETOACK(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDPMETOACK),
.CFGMSGRECEIVEDPMPME(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDPMPME),
.CFGMSGRECEIVEDSETSLOTPOWERLIMIT(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDSETSLOTPOWERLIMIT),
.CFGMSGRECEIVEDUNLOCK(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMSGRECEIVEDUNLOCK),
.CFGPCIECAPINTERRUPTMSGNUM({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CFGPCIELINKSTATE({PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIELINKSTATE2, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIELINKSTATE1, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIELINKSTATE0}),
.CFGPMCSRPMEEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMCSRPMEEN),
.CFGPMCSRPMESTATUS(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMCSRPMESTATUS),
.CFGPMCSRPOWERSTATE({PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMCSRPOWERSTATE1, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMCSRPOWERSTATE0}),
.CFGPMFORCESTATE({1'b0, 1'b0}),
.CFGPMFORCESTATEENN(1'b0),
.CFGPMHALTASPML0SN(1'b0),
.CFGPMHALTASPML1N(1'b0),
.CFGPMRCVASREQL1N(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMRCVASREQL1N),
.CFGPMRCVENTERL1N(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMRCVENTERL1N),
.CFGPMRCVENTERL23N(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMRCVENTERL23N),
.CFGPMRCVREQACKN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMRCVREQACKN),
.CFGPMSENDPMETON(1'b0),
.CFGPMTURNOFFOKN(1'b0),
.CFGPMWAKEN(1'b0),
.CFGPORTNUMBER({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CFGREVID({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CFGROOTCONTROLPMEINTEN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGROOTCONTROLPMEINTEN),
.CFGROOTCONTROLSYSERRCORRERREN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGROOTCONTROLSYSERRCORRERREN),
.CFGROOTCONTROLSYSERRFATALERREN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGROOTCONTROLSYSERRFATALERREN),
.CFGROOTCONTROLSYSERRNONFATALERREN(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGROOTCONTROLSYSERRNONFATALERREN),
.CFGSLOTCONTROLELECTROMECHILCTLPULSE(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSLOTCONTROLELECTROMECHILCTLPULSE),
.CFGSUBSYSID({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CFGSUBSYSVENDID({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CFGTRANSACTION(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTION),
.CFGTRANSACTIONADDR({PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONADDR6, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONADDR5, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONADDR4, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONADDR3, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONADDR2, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONADDR1, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONADDR0}),
.CFGTRANSACTIONTYPE(PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRANSACTIONTYPE),
.CFGTRNPENDINGN(1'b0),
.CFGVCTCVCMAP({PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVCTCVCMAP6, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVCTCVCMAP5, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVCTCVCMAP4, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVCTCVCMAP3, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVCTCVCMAP2, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVCTCVCMAP1, PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVCTCVCMAP0}),
.CFGVENDID({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.CMRSTN(1'b0),
.CMSTICKYRSTN(1'b0),
.DBGMODE({1'b0, 1'b0}),
.DBGSCLRA(PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRA),
.DBGSCLRB(PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRB),
.DBGSCLRC(PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRC),
.DBGSCLRD(PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRD),
.DBGSCLRE(PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRE),
.DBGSCLRF(PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRF),
.DBGSCLRG(PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRG),
.DBGSCLRH(PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRH),
.DBGSCLRI(PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRI),
.DBGSCLRJ(PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRJ),
.DBGSCLRK(PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSCLRK),
.DBGSUBMODE(1'b0),
.DBGVECA({PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA63, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA62, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA61, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA60, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA59, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA58, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA57, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA56, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA55, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA54, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA53, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA52, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA51, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA50, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA49, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA48, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA47, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA46, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA45, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA44, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA43, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA42, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA41, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA40, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA39, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA38, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA37, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA36, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA35, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA34, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA33, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA32, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA31, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA30, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA29, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA28, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA27, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA26, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA25, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA24, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA23, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA22, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA21, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA20, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA19, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA18, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA17, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA16, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA15, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA14, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA13, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA12, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA11, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA10, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA9, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA8, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA7, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA6, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA5, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA4, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA3, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA2, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA1, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECA0}),
.DBGVECB({PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB63, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB62, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB61, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB60, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB59, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB58, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB57, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB56, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB55, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB54, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB53, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB52, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB51, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB50, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB49, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB48, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB47, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB46, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB45, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB44, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB43, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB42, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB41, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB40, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB39, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB38, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB37, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB36, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB35, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB34, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB33, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB32, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB31, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB30, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB29, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB28, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB27, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB26, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB25, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB24, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB23, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB22, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB21, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB20, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB19, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB18, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB17, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB16, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB15, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB14, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB13, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB12, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB11, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB10, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB9, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB8, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB7, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB6, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB5, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB4, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB3, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB2, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB1, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECB0}),
.DBGVECC({PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC11, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC10, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC9, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC8, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC7, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC6, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC5, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC4, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC3, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC2, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC1, PCIE_BOT_X71Y115_PCIE_X0Y0_DBGVECC0}),
.DLRSTN(1'b0),
.DRPADDR({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.DRPCLK(1'b0),
.DRPDI({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.DRPDO({PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO15, PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO14, PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO13, PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO12, PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO11, PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO10, PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO9, PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO8, PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO7, PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO6, PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO5, PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO4, PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO3, PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO2, PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO1, PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDO0}),
.DRPEN(1'b0),
.DRPRDY(PCIE_BOT_X71Y115_PCIE_X0Y0_DRPRDY),
.DRPWE(1'b0),
.FUNCLVLRSTN(1'b0),
.LL2BADDLLPERR(PCIE_BOT_X71Y115_PCIE_X0Y0_LL2BADDLLPERR),
.LL2BADTLPERR(PCIE_BOT_X71Y115_PCIE_X0Y0_LL2BADTLPERR),
.LL2LINKSTATUS({PCIE_BOT_X71Y115_PCIE_X0Y0_LL2LINKSTATUS4, PCIE_BOT_X71Y115_PCIE_X0Y0_LL2LINKSTATUS3, PCIE_BOT_X71Y115_PCIE_X0Y0_LL2LINKSTATUS2, PCIE_BOT_X71Y115_PCIE_X0Y0_LL2LINKSTATUS1, PCIE_BOT_X71Y115_PCIE_X0Y0_LL2LINKSTATUS0}),
.LL2PROTOCOLERR(PCIE_BOT_X71Y115_PCIE_X0Y0_LL2PROTOCOLERR),
.LL2RECEIVERERR(PCIE_BOT_X71Y115_PCIE_X0Y0_LL2RECEIVERERR),
.LL2REPLAYROERR(PCIE_BOT_X71Y115_PCIE_X0Y0_LL2REPLAYROERR),
.LL2REPLAYTOERR(PCIE_BOT_X71Y115_PCIE_X0Y0_LL2REPLAYTOERR),
.LL2SENDASREQL1(1'b0),
.LL2SENDENTERL1(1'b0),
.LL2SENDENTERL23(1'b0),
.LL2SENDPMACK(1'b0),
.LL2SUSPENDNOW(1'b0),
.LL2SUSPENDOK(PCIE_BOT_X71Y115_PCIE_X0Y0_LL2SUSPENDOK),
.LL2TFCINIT1SEQ(PCIE_BOT_X71Y115_PCIE_X0Y0_LL2TFCINIT1SEQ),
.LL2TFCINIT2SEQ(PCIE_BOT_X71Y115_PCIE_X0Y0_LL2TFCINIT2SEQ),
.LL2TLPRCV(1'b0),
.LL2TXIDLE(PCIE_BOT_X71Y115_PCIE_X0Y0_LL2TXIDLE),
.LNKCLKEN(PCIE_BOT_X71Y115_PCIE_X0Y0_LNKCLKEN),
.MIMRXRADDR({PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR12, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR11, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR10, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR9, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR8, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR7, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR6, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR5, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR4, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR3, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR2, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR1, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRADDR0}),
.MIMRXRDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.MIMRXREN(PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXREN),
.MIMRXWADDR({PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR12, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR11, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR10, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR9, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR8, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR7, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR6, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR5, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR4, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR3, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR2, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR1, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWADDR0}),
.MIMRXWDATA({PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA67, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA66, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA65, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA64, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA63, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA62, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA61, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA60, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA59, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA58, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA57, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA56, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA55, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA54, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA53, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA52, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA51, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA50, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA49, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA48, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA47, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA46, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA45, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA44, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA43, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA42, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA41, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA40, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA39, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA38, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA37, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA36, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA35, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA34, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA33, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA32, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA31, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA30, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA29, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA28, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA27, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA26, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA25, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA24, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA23, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA22, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA21, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA20, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA19, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA18, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA17, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA16, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA15, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA14, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA13, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA12, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA11, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA10, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA9, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA8, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA7, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA6, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA5, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA4, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA3, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA2, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA1, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWDATA0}),
.MIMRXWEN(PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXWEN),
.MIMTXRADDR({PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR12, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR11, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR10, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR9, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR8, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR7, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR6, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR5, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR4, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR3, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR2, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR1, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRADDR0}),
.MIMTXRDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.MIMTXREN(PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXREN),
.MIMTXWADDR({PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR12, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR11, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR10, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR9, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR8, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR7, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR6, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR5, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR4, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR3, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR2, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR1, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWADDR0}),
.MIMTXWDATA({PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA68, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA67, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA66, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA65, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA64, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA63, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA62, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA61, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA60, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA59, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA58, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA57, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA56, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA55, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA54, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA53, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA52, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA51, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA50, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA49, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA48, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA47, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA46, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA45, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA44, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA43, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA42, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA41, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA40, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA39, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA38, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA37, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA36, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA35, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA34, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA33, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA32, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA31, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA30, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA29, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA28, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA27, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA26, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA25, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA24, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA23, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA22, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA21, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA20, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA19, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA18, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA17, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA16, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA15, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA14, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA13, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA12, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA11, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA10, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA9, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA8, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA7, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA6, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA5, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA4, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA3, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA2, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA1, PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWDATA0}),
.MIMTXWEN(PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXWEN),
.PIPECLK(1'b0),
.PIPERX0CHANISALIGNED(1'b0),
.PIPERX0CHARISK({1'b0, 1'b0}),
.PIPERX0DATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.PIPERX0ELECIDLE(1'b0),
.PIPERX0PHYSTATUS(1'b0),
.PIPERX0POLARITY(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0POLARITY),
.PIPERX0STATUS({1'b0, 1'b0, 1'b0}),
.PIPERX0VALID(1'b0),
.PIPERX1CHANISALIGNED(1'b0),
.PIPERX1CHARISK({1'b0, 1'b0}),
.PIPERX1DATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.PIPERX1ELECIDLE(1'b0),
.PIPERX1PHYSTATUS(1'b0),
.PIPERX1POLARITY(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1POLARITY),
.PIPERX1STATUS({1'b0, 1'b0, 1'b0}),
.PIPERX1VALID(1'b0),
.PIPERX2CHANISALIGNED(1'b0),
.PIPERX2CHARISK({1'b0, 1'b0}),
.PIPERX2DATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.PIPERX2ELECIDLE(1'b0),
.PIPERX2PHYSTATUS(1'b0),
.PIPERX2POLARITY(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2POLARITY),
.PIPERX2STATUS({1'b0, 1'b0, 1'b0}),
.PIPERX2VALID(1'b0),
.PIPERX3CHANISALIGNED(1'b0),
.PIPERX3CHARISK({1'b0, 1'b0}),
.PIPERX3DATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.PIPERX3ELECIDLE(1'b0),
.PIPERX3PHYSTATUS(1'b0),
.PIPERX3POLARITY(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3POLARITY),
.PIPERX3STATUS({1'b0, 1'b0, 1'b0}),
.PIPERX3VALID(1'b0),
.PIPERX4CHANISALIGNED(1'b0),
.PIPERX4CHARISK({1'b0, 1'b0}),
.PIPERX4DATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.PIPERX4ELECIDLE(1'b0),
.PIPERX4PHYSTATUS(1'b0),
.PIPERX4POLARITY(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4POLARITY),
.PIPERX4STATUS({1'b0, 1'b0, 1'b0}),
.PIPERX4VALID(1'b0),
.PIPERX5CHANISALIGNED(1'b0),
.PIPERX5CHARISK({1'b0, 1'b0}),
.PIPERX5DATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.PIPERX5ELECIDLE(1'b0),
.PIPERX5PHYSTATUS(1'b0),
.PIPERX5POLARITY(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5POLARITY),
.PIPERX5STATUS({1'b0, 1'b0, 1'b0}),
.PIPERX5VALID(1'b0),
.PIPERX6CHANISALIGNED(1'b0),
.PIPERX6CHARISK({1'b0, 1'b0}),
.PIPERX6DATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.PIPERX6ELECIDLE(1'b0),
.PIPERX6PHYSTATUS(1'b0),
.PIPERX6POLARITY(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6POLARITY),
.PIPERX6STATUS({1'b0, 1'b0, 1'b0}),
.PIPERX6VALID(1'b0),
.PIPERX7CHANISALIGNED(1'b0),
.PIPERX7CHARISK({1'b0, 1'b0}),
.PIPERX7DATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.PIPERX7ELECIDLE(1'b0),
.PIPERX7PHYSTATUS(1'b0),
.PIPERX7POLARITY(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7POLARITY),
.PIPERX7STATUS({1'b0, 1'b0, 1'b0}),
.PIPERX7VALID(1'b0),
.PIPETX0CHARISK({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0CHARISK1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0CHARISK0}),
.PIPETX0COMPLIANCE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0COMPLIANCE),
.PIPETX0DATA({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA15, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA14, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA13, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA12, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA11, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA10, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA9, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA8, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA7, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA6, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA5, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA4, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA3, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA2, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0DATA0}),
.PIPETX0ELECIDLE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0ELECIDLE),
.PIPETX0POWERDOWN({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0POWERDOWN1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX0POWERDOWN0}),
.PIPETX1CHARISK({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1CHARISK1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1CHARISK0}),
.PIPETX1COMPLIANCE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1COMPLIANCE),
.PIPETX1DATA({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA15, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA14, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA13, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA12, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA11, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA10, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA9, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA8, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA7, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA6, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA5, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA4, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA3, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA2, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1DATA0}),
.PIPETX1ELECIDLE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1ELECIDLE),
.PIPETX1POWERDOWN({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1POWERDOWN1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX1POWERDOWN0}),
.PIPETX2CHARISK({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2CHARISK1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2CHARISK0}),
.PIPETX2COMPLIANCE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2COMPLIANCE),
.PIPETX2DATA({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA15, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA14, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA13, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA12, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA11, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA10, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA9, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA8, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA7, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA6, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA5, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA4, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA3, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA2, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2DATA0}),
.PIPETX2ELECIDLE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2ELECIDLE),
.PIPETX2POWERDOWN({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2POWERDOWN1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX2POWERDOWN0}),
.PIPETX3CHARISK({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3CHARISK1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3CHARISK0}),
.PIPETX3COMPLIANCE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3COMPLIANCE),
.PIPETX3DATA({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA15, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA14, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA13, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA12, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA11, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA10, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA9, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA8, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA7, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA6, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA5, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA4, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA3, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA2, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3DATA0}),
.PIPETX3ELECIDLE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3ELECIDLE),
.PIPETX3POWERDOWN({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3POWERDOWN1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX3POWERDOWN0}),
.PIPETX4CHARISK({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4CHARISK1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4CHARISK0}),
.PIPETX4COMPLIANCE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4COMPLIANCE),
.PIPETX4DATA({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA15, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA14, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA13, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA12, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA11, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA10, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA9, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA8, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA7, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA6, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA5, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA4, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA3, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA2, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4DATA0}),
.PIPETX4ELECIDLE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4ELECIDLE),
.PIPETX4POWERDOWN({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4POWERDOWN1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX4POWERDOWN0}),
.PIPETX5CHARISK({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5CHARISK1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5CHARISK0}),
.PIPETX5COMPLIANCE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5COMPLIANCE),
.PIPETX5DATA({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA15, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA14, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA13, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA12, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA11, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA10, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA9, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA8, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA7, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA6, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA5, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA4, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA3, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA2, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5DATA0}),
.PIPETX5ELECIDLE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5ELECIDLE),
.PIPETX5POWERDOWN({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5POWERDOWN1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX5POWERDOWN0}),
.PIPETX6CHARISK({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6CHARISK1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6CHARISK0}),
.PIPETX6COMPLIANCE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6COMPLIANCE),
.PIPETX6DATA({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA15, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA14, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA13, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA12, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA11, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA10, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA9, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA8, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA7, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA6, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA5, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA4, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA3, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA2, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6DATA0}),
.PIPETX6ELECIDLE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6ELECIDLE),
.PIPETX6POWERDOWN({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6POWERDOWN1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX6POWERDOWN0}),
.PIPETX7CHARISK({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7CHARISK1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7CHARISK0}),
.PIPETX7COMPLIANCE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7COMPLIANCE),
.PIPETX7DATA({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA15, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA14, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA13, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA12, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA11, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA10, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA9, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA8, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA7, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA6, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA5, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA4, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA3, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA2, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7DATA0}),
.PIPETX7ELECIDLE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7ELECIDLE),
.PIPETX7POWERDOWN({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7POWERDOWN1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETX7POWERDOWN0}),
.PIPETXDEEMPH(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETXDEEMPH),
.PIPETXMARGIN({PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETXMARGIN2, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETXMARGIN1, PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETXMARGIN0}),
.PIPETXRATE(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETXRATE),
.PIPETXRCVRDET(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETXRCVRDET),
.PIPETXRESET(PCIE_BOT_X71Y115_PCIE_X0Y0_PIPETXRESET),
.PL2DIRECTEDLSTATE({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.PL2L0REQ(PCIE_BOT_X71Y115_PCIE_X0Y0_PL2L0REQ),
.PL2LINKUP(PCIE_BOT_X71Y115_PCIE_X0Y0_PL2LINKUP),
.PL2RECEIVERERR(PCIE_BOT_X71Y115_PCIE_X0Y0_PL2RECEIVERERR),
.PL2RECOVERY(PCIE_BOT_X71Y115_PCIE_X0Y0_PL2RECOVERY),
.PL2RXELECIDLE(PCIE_BOT_X71Y115_PCIE_X0Y0_PL2RXELECIDLE),
.PL2RXPMSTATE({PCIE_BOT_X71Y115_PCIE_X0Y0_PL2RXPMSTATE1, PCIE_BOT_X71Y115_PCIE_X0Y0_PL2RXPMSTATE0}),
.PL2SUSPENDOK(PCIE_BOT_X71Y115_PCIE_X0Y0_PL2SUSPENDOK),
.PLDBGMODE({1'b0, 1'b0, 1'b0}),
.PLDBGVEC({PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC11, PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC10, PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC9, PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC8, PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC7, PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC6, PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC5, PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC4, PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC3, PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC2, PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC1, PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGVEC0}),
.PLDIRECTEDCHANGEDONE(PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDCHANGEDONE),
.PLDIRECTEDLINKAUTON(1'b0),
.PLDIRECTEDLINKCHANGE({1'b0, 1'b0}),
.PLDIRECTEDLINKSPEED(1'b0),
.PLDIRECTEDLINKWIDTH({1'b0, 1'b0}),
.PLDIRECTEDLTSSMNEW({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.PLDIRECTEDLTSSMNEWVLD(1'b0),
.PLDIRECTEDLTSSMSTALL(1'b0),
.PLDOWNSTREAMDEEMPHSOURCE(1'b0),
.PLINITIALLINKWIDTH({PCIE_BOT_X71Y115_PCIE_X0Y0_PLINITIALLINKWIDTH2, PCIE_BOT_X71Y115_PCIE_X0Y0_PLINITIALLINKWIDTH1, PCIE_BOT_X71Y115_PCIE_X0Y0_PLINITIALLINKWIDTH0}),
.PLLANEREVERSALMODE({PCIE_BOT_X71Y115_PCIE_X0Y0_PLLANEREVERSALMODE1, PCIE_BOT_X71Y115_PCIE_X0Y0_PLLANEREVERSALMODE0}),
.PLLINKGEN2CAP(PCIE_BOT_X71Y115_PCIE_X0Y0_PLLINKGEN2CAP),
.PLLINKPARTNERGEN2SUPPORTED(PCIE_BOT_X71Y115_PCIE_X0Y0_PLLINKPARTNERGEN2SUPPORTED),
.PLLINKUPCFGCAP(PCIE_BOT_X71Y115_PCIE_X0Y0_PLLINKUPCFGCAP),
.PLLTSSMSTATE({PCIE_BOT_X71Y115_PCIE_X0Y0_PLLTSSMSTATE5, PCIE_BOT_X71Y115_PCIE_X0Y0_PLLTSSMSTATE4, PCIE_BOT_X71Y115_PCIE_X0Y0_PLLTSSMSTATE3, PCIE_BOT_X71Y115_PCIE_X0Y0_PLLTSSMSTATE2, PCIE_BOT_X71Y115_PCIE_X0Y0_PLLTSSMSTATE1, PCIE_BOT_X71Y115_PCIE_X0Y0_PLLTSSMSTATE0}),
.PLPHYLNKUPN(PCIE_BOT_X71Y115_PCIE_X0Y0_PLPHYLNKUPN),
.PLRECEIVEDHOTRST(PCIE_BOT_X71Y115_PCIE_X0Y0_PLRECEIVEDHOTRST),
.PLRSTN(1'b0),
.PLRXPMSTATE({PCIE_BOT_X71Y115_PCIE_X0Y0_PLRXPMSTATE1, PCIE_BOT_X71Y115_PCIE_X0Y0_PLRXPMSTATE0}),
.PLSELLNKRATE(PCIE_BOT_X71Y115_PCIE_X0Y0_PLSELLNKRATE),
.PLSELLNKWIDTH({PCIE_BOT_X71Y115_PCIE_X0Y0_PLSELLNKWIDTH1, PCIE_BOT_X71Y115_PCIE_X0Y0_PLSELLNKWIDTH0}),
.PLTRANSMITHOTRST(1'b0),
.PLTXPMSTATE({PCIE_BOT_X71Y115_PCIE_X0Y0_PLTXPMSTATE2, PCIE_BOT_X71Y115_PCIE_X0Y0_PLTXPMSTATE1, PCIE_BOT_X71Y115_PCIE_X0Y0_PLTXPMSTATE0}),
.PLUPSTREAMPREFERDEEMPH(1'b0),
.RECEIVEDFUNCLVLRSTN(PCIE_BOT_X71Y115_PCIE_X0Y0_RECEIVEDFUNCLVLRSTN),
.SYSRSTN(LIOB33_X0Y11_IOB_X0Y11_I),
.TL2ASPMSUSPENDCREDITCHECK(1'b0),
.TL2ASPMSUSPENDCREDITCHECKOK(PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ASPMSUSPENDCREDITCHECKOK),
.TL2ASPMSUSPENDREQ(PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ASPMSUSPENDREQ),
.TL2ERRFCPE(PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRFCPE),
.TL2ERRHDR({PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR63, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR62, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR61, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR60, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR59, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR58, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR57, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR56, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR55, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR54, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR53, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR52, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR51, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR50, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR49, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR48, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR47, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR46, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR45, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR44, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR43, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR42, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR41, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR40, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR39, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR38, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR37, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR36, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR35, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR34, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR33, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR32, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR31, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR30, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR29, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR28, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR27, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR26, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR25, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR24, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR23, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR22, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR21, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR20, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR19, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR18, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR17, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR16, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR15, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR14, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR13, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR12, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR11, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR10, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR9, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR8, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR7, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR6, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR5, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR4, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR3, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR2, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR1, PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRHDR0}),
.TL2ERRMALFORMED(PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRMALFORMED),
.TL2ERRRXOVERFLOW(PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ERRRXOVERFLOW),
.TL2PPMSUSPENDOK(PCIE_BOT_X71Y115_PCIE_X0Y0_TL2PPMSUSPENDOK),
.TL2PPMSUSPENDREQ(1'b0),
.TLRSTN(1'b0),
.TRNFCCPLD({PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD11, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD10, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD9, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD8, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD7, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD6, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD5, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD4, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD3, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD2, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD1, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLD0}),
.TRNFCCPLH({PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH7, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH6, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH5, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH4, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH3, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH2, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH1, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCCPLH0}),
.TRNFCNPD({PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD11, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD10, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD9, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD8, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD7, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD6, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD5, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD4, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD3, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD2, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD1, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPD0}),
.TRNFCNPH({PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH7, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH6, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH5, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH4, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH3, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH2, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH1, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCNPH0}),
.TRNFCPD({PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD11, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD10, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD9, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD8, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD7, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD6, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD5, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD4, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD3, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD2, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD1, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPD0}),
.TRNFCPH({PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH7, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH6, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH5, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH4, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH3, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH2, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH1, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCPH0}),
.TRNFCSEL({1'b0, 1'b0, 1'b0}),
.TRNLNKUP(PCIE_BOT_X71Y115_PCIE_X0Y0_TRNLNKUP),
.TRNRBARHIT({PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT7, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT6, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT5, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT4, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT3, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT2, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT1, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRBARHIT0}),
.TRNRD({PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD127, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD126, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD125, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD124, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD123, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD122, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD121, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD120, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD119, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD118, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD117, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD116, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD115, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD114, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD113, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD112, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD111, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD110, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD109, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD108, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD107, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD106, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD105, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD104, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD103, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD102, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD101, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD100, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD99, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD98, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD97, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD96, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD95, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD94, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD93, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD92, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD91, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD90, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD89, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD88, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD87, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD86, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD85, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD84, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD83, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD82, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD81, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD80, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD79, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD78, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD77, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD76, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD75, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD74, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD73, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD72, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD71, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD70, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD69, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD68, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD67, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD66, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD65, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD64, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD63, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD62, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD61, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD60, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD59, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD58, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD57, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD56, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD55, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD54, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD53, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD52, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD51, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD50, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD49, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD48, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD47, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD46, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD45, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD44, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD43, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD42, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD41, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD40, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD39, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD38, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD37, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD36, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD35, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD34, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD33, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD32, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD31, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD30, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD29, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD28, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD27, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD26, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD25, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD24, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD23, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD22, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD21, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD20, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD19, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD18, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD17, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD16, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD15, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD14, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD13, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD12, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD11, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD10, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD9, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD8, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD7, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD6, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD5, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD4, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD3, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD2, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD1, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRD0}),
.TRNRDLLPDATA({PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA63, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA62, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA61, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA60, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA59, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA58, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA57, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA56, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA55, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA54, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA53, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA52, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA51, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA50, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA49, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA48, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA47, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA46, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA45, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA44, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA43, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA42, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA41, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA40, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA39, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA38, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA37, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA36, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA35, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA34, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA33, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA32, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA31, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA30, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA29, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA28, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA27, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA26, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA25, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA24, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA23, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA22, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA21, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA20, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA19, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA18, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA17, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA16, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA15, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA14, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA13, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA12, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA11, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA10, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA9, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA8, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA7, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA6, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA5, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA4, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA3, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA2, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA1, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPDATA0}),
.TRNRDLLPSRCRDY({PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPSRCRDY1, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDLLPSRCRDY0}),
.TRNRDSTRDY(1'b0),
.TRNRECRCERR(PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRECRCERR),
.TRNREOF(PCIE_BOT_X71Y115_PCIE_X0Y0_TRNREOF),
.TRNRERRFWD(PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRERRFWD),
.TRNRFCPRET(1'b0),
.TRNRNPOK(1'b0),
.TRNRNPREQ(1'b0),
.TRNRREM({PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRREM1, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRREM0}),
.TRNRSOF(PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRSOF),
.TRNRSRCDSC(PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRSRCDSC),
.TRNRSRCRDY(PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRSRCRDY),
.TRNTBUFAV({PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTBUFAV5, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTBUFAV4, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTBUFAV3, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTBUFAV2, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTBUFAV1, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTBUFAV0}),
.TRNTCFGGNT(1'b0),
.TRNTCFGREQ(PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTCFGREQ),
.TRNTD({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.TRNTDLLPDATA({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}),
.TRNTDLLPDSTRDY(PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDSTRDY),
.TRNTDLLPSRCRDY(1'b0),
.TRNTDSTRDY({PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDSTRDY3, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDSTRDY2, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDSTRDY1, PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDSTRDY0}),
.TRNTECRCGEN(1'b0),
.TRNTEOF(1'b0),
.TRNTERRDROP(PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTERRDROP),
.TRNTERRFWD(1'b0),
.TRNTREM({1'b0, 1'b0}),
.TRNTSOF(1'b0),
.TRNTSRCDSC(1'b0),
.TRNTSRCRDY(1'b0),
.TRNTSTR(1'b0),
.USERCLK(1'b0),
.USERCLK2(1'b0),
.USERRSTN(PCIE_BOT_X71Y115_PCIE_X0Y0_USERRSTN)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y31_IOB_X1Y32_OBUF (
.I(RIOB33_X43Y45_IOB_X1Y46_I),
.O(led[11])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y37_IOB_X1Y37_OBUF (
.I(RIOB33_X43Y47_IOB_X1Y47_I),
.O(led[10])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y37_IOB_X1Y38_OBUF (
.I(RIOB33_X43Y45_IOB_X1Y45_I),
.O(led[9])
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y39_IOB_X1Y39_IBUF (
.I(sw[12]),
.O(RIOB33_X43Y39_IOB_X1Y39_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y39_IOB_X1Y40_IBUF (
.I(sw[8]),
.O(RIOB33_X43Y39_IOB_X1Y40_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y43_IOB_X1Y43_IBUF (
.I(sw[13]),
.O(RIOB33_X43Y43_IOB_X1Y43_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y43_IOB_X1Y44_IBUF (
.I(sw[14]),
.O(RIOB33_X43Y43_IOB_X1Y44_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y45_IOB_X1Y45_IBUF (
.I(sw[9]),
.O(RIOB33_X43Y45_IOB_X1Y45_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y45_IOB_X1Y46_IBUF (
.I(sw[11]),
.O(RIOB33_X43Y45_IOB_X1Y46_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y47_IOB_X1Y47_IBUF (
.I(sw[10]),
.O(RIOB33_X43Y47_IOB_X1Y47_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) RIOB33_X43Y47_IOB_X1Y48_IBUF (
.I(sw[15]),
.O(RIOB33_X43Y47_IOB_X1Y48_I)
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y61_IOB_X1Y61_OBUF (
.I(RIOB33_X43Y43_IOB_X1Y44_I),
.O(led[14])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y75_IOB_X1Y75_OBUF (
.I(RIOB33_X43Y39_IOB_X1Y39_I),
.O(led[12])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y75_IOB_X1Y76_OBUF (
.I(RIOB33_X43Y43_IOB_X1Y43_I),
.O(led[13])
  );


  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) RIOB33_X43Y87_IOB_X1Y87_OBUF (
.I(RIOB33_X43Y47_IOB_X1Y48_I),
.O(led[15])
  );
  assign LIOI3_X0Y1_OLOGIC_X0Y2_OQ = RIOB33_X43Y39_IOB_X1Y40_I;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_TQ = 1'b1;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_OQ = LIOB33_X0Y5_IOB_X0Y6_I;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_TQ = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_OQ = LIOB33_X0Y7_IOB_X0Y8_I;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_TQ = 1'b1;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_OQ = PCIE_BOT_X71Y115_PCIE_X0Y0_DRPRDY;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_TQ = 1'b1;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_O = LIOB33_X0Y5_IOB_X0Y6_I;
  assign LIOI3_X0Y5_ILOGIC_X0Y5_O = LIOB33_X0Y5_IOB_X0Y5_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_O = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y9_O = LIOB33_X0Y9_IOB_X0Y9_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_O = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_O = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_OQ = LIOB33_X0Y7_IOB_X0Y7_I;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_TQ = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_OQ = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_TQ = 1'b1;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_OQ = LIOB33_X0Y5_IOB_X0Y5_I;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_O = LIOB33_X0Y7_IOB_X0Y8_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_O = LIOB33_X0Y7_IOB_X0Y7_I;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_OQ = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_OQ = LIOB33_X0Y9_IOB_X0Y9_I;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ = 1'b1;
  assign RIOI3_X43Y39_ILOGIC_X1Y40_O = RIOB33_X43Y39_IOB_X1Y40_I;
  assign RIOI3_X43Y39_ILOGIC_X1Y39_O = RIOB33_X43Y39_IOB_X1Y39_I;
  assign RIOI3_X43Y45_ILOGIC_X1Y46_O = RIOB33_X43Y45_IOB_X1Y46_I;
  assign RIOI3_X43Y45_ILOGIC_X1Y45_O = RIOB33_X43Y45_IOB_X1Y45_I;
  assign RIOI3_X43Y47_ILOGIC_X1Y48_O = RIOB33_X43Y47_IOB_X1Y48_I;
  assign RIOI3_X43Y47_ILOGIC_X1Y47_O = RIOB33_X43Y47_IOB_X1Y47_I;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_OQ = RIOB33_X43Y43_IOB_X1Y44_I;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_TQ = 1'b1;
  assign RIOI3_X43Y75_OLOGIC_X1Y76_OQ = RIOB33_X43Y43_IOB_X1Y43_I;
  assign RIOI3_X43Y75_OLOGIC_X1Y76_TQ = 1'b1;
  assign RIOI3_X43Y75_OLOGIC_X1Y75_OQ = RIOB33_X43Y39_IOB_X1Y39_I;
  assign RIOI3_X43Y75_OLOGIC_X1Y75_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_OQ = RIOB33_X43Y45_IOB_X1Y46_I;
  assign RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_TQ = 1'b1;
  assign RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_O = RIOB33_X43Y43_IOB_X1Y44_I;
  assign RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_O = RIOB33_X43Y43_IOB_X1Y43_I;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_OQ = RIOB33_X43Y45_IOB_X1Y45_I;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_OQ = RIOB33_X43Y47_IOB_X1Y47_I;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_TQ = 1'b1;
  assign RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_OQ = RIOB33_X43Y47_IOB_X1Y48_I;
  assign RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_TQ = 1'b1;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPECLK = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0CHANISALIGNED = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0CHARISK0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0CHARISK1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0DATA15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0ELECIDLE = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0PHYSTATUS = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0STATUS0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0STATUS1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0STATUS2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX0VALID = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1CHANISALIGNED = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1CHARISK0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1CHARISK1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1DATA15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1ELECIDLE = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1PHYSTATUS = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1STATUS0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1STATUS1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1STATUS2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX1VALID = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2CHANISALIGNED = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2CHARISK0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2CHARISK1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2DATA15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2ELECIDLE = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2PHYSTATUS = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2STATUS0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2STATUS1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2STATUS2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX2VALID = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3CHANISALIGNED = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3CHARISK0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3CHARISK1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3DATA15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3ELECIDLE = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3PHYSTATUS = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3STATUS0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3STATUS1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_FUNCLVLRSTN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3STATUS2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX3VALID = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4CHANISALIGNED = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4CHARISK0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4CHARISK1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4DATA15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4ELECIDLE = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4PHYSTATUS = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4STATUS0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4STATUS1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4STATUS2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX4VALID = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5CHANISALIGNED = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5CHARISK0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5CHARISK1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA13 = 1'b0;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_D = LIOB33_X0Y5_IOB_X0Y6_I;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5DATA15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5ELECIDLE = 1'b0;
  assign LIOI3_X0Y5_ILOGIC_X0Y5_D = LIOB33_X0Y5_IOB_X0Y5_I;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5PHYSTATUS = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5STATUS0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5STATUS1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5STATUS2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX5VALID = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6CHANISALIGNED = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6CHARISK0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6CHARISK1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6DATA15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6ELECIDLE = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6PHYSTATUS = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6STATUS0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6STATUS1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6STATUS2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX6VALID = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7CHANISALIGNED = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7CHARISK0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7CHARISK1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7DATA15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7ELECIDLE = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7PHYSTATUS = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7STATUS0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7STATUS1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7STATUS2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PIPERX7VALID = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PL2DIRECTEDLSTATE0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PL2DIRECTEDLSTATE1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PL2DIRECTEDLSTATE2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PL2DIRECTEDLSTATE3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PL2DIRECTEDLSTATE4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGMODE0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGMODE1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDBGMODE2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLINKAUTON = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLINKCHANGE0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLINKCHANGE1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLINKSPEED = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLINKWIDTH0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLINKWIDTH1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMNEW0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMNEW1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMNEW2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMNEW3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMNEW4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMNEW5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMNEWVLD = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDIRECTEDLTSSMSTALL = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLDOWNSTREAMDEEMPHSOURCE = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLRSTN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLTRANSMITHOTRST = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_PLUPSTREAMPREFERDEEMPH = 1'b0;
  assign LIOB33_X0Y43_IOB_X0Y43_O = LIOB33_X0Y11_IOB_X0Y12_I;
  assign RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_D1 = RIOB33_X43Y47_IOB_X1Y48_I;
  assign RIOI3_TBYTETERM_X43Y87_OLOGIC_X1Y87_T1 = 1'b1;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_D = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y9_D = LIOB33_X0Y9_IOB_X0Y9_I;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_D1 = RIOB33_X43Y43_IOB_X1Y44_I;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_SYSRSTN = LIOB33_X0Y11_IOB_X0Y11_I;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TL2ASPMSUSPENDCREDITCHECK = 1'b0;
  assign RIOI3_X43Y61_OLOGIC_X1Y61_T1 = 1'b1;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TL2PPMSUSPENDREQ = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TLRSTN = 1'b0;
  assign RIOI3_X43Y75_OLOGIC_X1Y76_D1 = RIOB33_X43Y43_IOB_X1Y43_I;
  assign RIOI3_X43Y75_OLOGIC_X1Y76_T1 = 1'b1;
  assign RIOI3_X43Y75_OLOGIC_X1Y75_D1 = RIOB33_X43Y39_IOB_X1Y39_I;
  assign RIOI3_X43Y75_OLOGIC_X1Y75_T1 = 1'b1;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCSEL0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCSEL1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNFCSEL2 = 1'b0;
  assign LIOB33_X0Y17_IOB_X0Y18_O = LIOB33_X0Y7_IOB_X0Y7_I;
  assign RIOB33_X43Y87_IOB_X1Y87_O = RIOB33_X43Y47_IOB_X1Y48_I;
  assign RIOI3_X43Y45_ILOGIC_X1Y46_D = RIOB33_X43Y45_IOB_X1Y46_I;
  assign RIOI3_X43Y45_ILOGIC_X1Y45_D = RIOB33_X43Y45_IOB_X1Y45_I;
  assign RIOB33_X43Y37_IOB_X1Y38_O = RIOB33_X43Y45_IOB_X1Y45_I;
  assign RIOB33_X43Y37_IOB_X1Y37_O = RIOB33_X43Y47_IOB_X1Y47_I;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRDSTRDY = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRFCPRET = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRNPOK = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNRNPREQ = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTCFGGNT = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD16 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD17 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD18 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD19 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD20 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD21 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD22 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD23 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD24 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD25 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD26 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD27 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD28 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD29 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD30 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD31 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD32 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD33 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD34 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD35 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD36 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD37 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD38 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD39 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD40 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD41 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD42 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD43 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD44 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD45 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD46 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD47 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD48 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD49 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD50 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD51 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD52 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD53 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD54 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD55 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD56 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD57 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD58 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD59 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD60 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD61 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD62 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD63 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD64 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD65 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD66 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD67 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD68 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD69 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD70 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD71 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD72 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD73 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD74 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD75 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD76 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD77 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD78 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD79 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD80 = 1'b0;
  assign LIOB33_X0Y19_IOB_X0Y20_O = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOB33_X0Y19_IOB_X0Y19_O = LIOB33_X0Y9_IOB_X0Y9_I;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD81 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD82 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD83 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD84 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD85 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD86 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD87 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD88 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD89 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD90 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD91 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD92 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD93 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD94 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD95 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD96 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD97 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD98 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD99 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD100 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD101 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD102 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD103 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD104 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD105 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD106 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD107 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD108 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD109 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD110 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD111 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD112 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD113 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD114 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD115 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD116 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD117 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD118 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD119 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD120 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD121 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD122 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD123 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD124 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD125 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD126 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTD127 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA16 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA17 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA18 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA19 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA20 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA21 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA22 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA23 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA24 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA25 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA26 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA27 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA28 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA29 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA30 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPDATA31 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTDLLPSRCRDY = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTECRCGEN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTEOF = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTERRFWD = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTREM0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTREM1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTSOF = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTSRCDSC = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTSRCRDY = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_TRNTSTR = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_USERCLK = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_USERCLK2 = 1'b0;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_T1 = 1'b1;
  assign RIOB33_X43Y61_IOB_X1Y61_O = RIOB33_X43Y43_IOB_X1Y44_I;
  assign LIOB33_X0Y111_IOB_X0Y111_O = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_D = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_D = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_D = LIOB33_X0Y7_IOB_X0Y8_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_D = LIOB33_X0Y7_IOB_X0Y7_I;
  assign RIOB33_X43Y31_IOB_X1Y32_O = RIOB33_X43Y45_IOB_X1Y46_I;
  assign RIOI3_X43Y47_ILOGIC_X1Y48_D = RIOB33_X43Y47_IOB_X1Y48_I;
  assign RIOI3_X43Y47_ILOGIC_X1Y47_D = RIOB33_X43Y47_IOB_X1Y47_I;
  assign LIOB33_SING_X0Y0_IOB_X0Y0_O = LIOB33_X0Y5_IOB_X0Y5_I;
  assign RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_D1 = RIOB33_X43Y45_IOB_X1Y46_I;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_D1 = LIOB33_X0Y9_IOB_X0Y10_I;
  assign RIOI3_TBYTESRC_X43Y31_OLOGIC_X1Y32_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y20_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_D1 = LIOB33_X0Y9_IOB_X0Y9_I;
  assign LIOI3_TBYTESRC_X0Y19_OLOGIC_X0Y19_T1 = 1'b1;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERINTERRUPTMSGNUM0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERINTERRUPTMSGNUM1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERINTERRUPTMSGNUM2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERINTERRUPTMSGNUM3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGAERINTERRUPTMSGNUM4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_LL2SENDASREQL1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_LL2SENDENTERL1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_LL2SENDENTERL23 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_LL2SENDPMACK = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_LL2SUSPENDNOW = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDEVID15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSBUSNUMBER7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSDEVICENUMBER0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSDEVICENUMBER1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSDEVICENUMBER2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSDEVICENUMBER3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSDEVICENUMBER4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSFUNCTIONNUMBER0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSFUNCTIONNUMBER1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSFUNCTIONNUMBER2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN16 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN17 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN18 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN19 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN20 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN21 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN22 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN23 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN24 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN25 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN26 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN27 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN28 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN29 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN30 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN31 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN32 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN33 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN34 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN35 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN36 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN37 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN38 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN39 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN40 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN41 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN42 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN43 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN44 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN45 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN46 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN47 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN48 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN49 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN50 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN51 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN52 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN53 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN54 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN55 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN56 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN57 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN58 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN59 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN60 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN61 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN62 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGDSN63 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRACSN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG16 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG17 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG18 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG19 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG20 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG21 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG22 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG23 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG24 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG25 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG26 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG27 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG28 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG29 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG30 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG31 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG32 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG33 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG34 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG35 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG36 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG37 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG38 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG39 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG40 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG41 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG42 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG43 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG44 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG45 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG46 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG47 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG48 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG49 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG50 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG51 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG52 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG53 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG54 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG55 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG56 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG57 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG58 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG59 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG60 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG61 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG62 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG63 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG64 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG65 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG66 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG67 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG68 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG69 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG70 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG71 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG72 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG73 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG74 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG75 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG76 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG77 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG78 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG79 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG80 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG81 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG82 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG83 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG84 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG85 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG86 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG87 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG88 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG89 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG90 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG91 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG92 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG93 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG94 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG95 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG96 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG97 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG98 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG99 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG100 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG101 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG102 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG103 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG104 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG105 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG106 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG107 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG108 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG109 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG110 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG111 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG112 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG113 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG114 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG115 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG116 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG117 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG118 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG119 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG120 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG121 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG122 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG123 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG124 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG125 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG126 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRAERHEADERLOG127 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRATOMICEGRESSBLOCKEDN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRCORN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRCPLABORTN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRCPLTIMEOUTN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRCPLUNEXPECTN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRECRCN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRINTERNALCORN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRINTERNALUNCORN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRLOCKEDN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRMALFORMEDN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRMCBLOCKEDN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRNORECOVERYN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRPOISONEDN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRPOSTEDN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER16 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER17 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER18 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER19 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER20 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER21 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER22 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER23 = 1'b0;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_D1 = RIOB33_X43Y39_IOB_X1Y40_I;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER24 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER25 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER26 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER27 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER28 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER29 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER30 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER31 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER32 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER33 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER34 = 1'b0;
  assign LIOI3_X0Y1_OLOGIC_X0Y2_T1 = 1'b1;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER35 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER36 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER37 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER38 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER39 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER40 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER41 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER42 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER43 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER44 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER45 = 1'b0;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_D1 = LIOB33_X0Y5_IOB_X0Y6_I;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER46 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRTLPCPLHEADER47 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGERRURN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGFORCECOMMONCLOCKOFF = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGFORCEEXTENDEDSYNCON = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGFORCEMPS0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGFORCEMPS1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGFORCEMPS2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTASSERTN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI1 = 1'b0;
  assign LIOI3_X0Y1_OLOGIC_X0Y1_T1 = 1'b1;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTDI7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGINTERRUPTSTATN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTBYTEENN0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTBYTEENN1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTBYTEENN2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTBYTEENN3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI16 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI17 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI18 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI19 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI20 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI21 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI22 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI23 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI24 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI25 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI26 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI27 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI28 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI29 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI30 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDI31 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTDWADDR9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTRDENN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTWRENN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTWRREADONLYN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGMGMTWRRW1CASRWN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIECAPINTERRUPTMSGNUM0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIECAPINTERRUPTMSGNUM1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIECAPINTERRUPTMSGNUM2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIECAPINTERRUPTMSGNUM3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPCIECAPINTERRUPTMSGNUM4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMFORCESTATE0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMFORCESTATE1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMFORCESTATEENN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMHALTASPML0SN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMHALTASPML1N = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMSENDPMETON = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMTURNOFFOKN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPMWAKEN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGPORTNUMBER7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGREVID7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSID15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGSUBSYSVENDID15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGTRNPENDINGN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CFGVENDID15 = 1'b0;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_D1 = LIOB33_X0Y7_IOB_X0Y7_I;
  assign LIOI3_X0Y17_OLOGIC_X0Y18_T1 = 1'b1;
  assign LIOB33_X0Y1_IOB_X0Y2_O = RIOB33_X43Y39_IOB_X1Y40_I;
  assign LIOB33_X0Y1_IOB_X0Y1_O = LIOB33_X0Y5_IOB_X0Y6_I;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CMRSTN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_CMSTICKYRSTN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DBGMODE0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DBGMODE1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DBGSUBMODE = 1'b0;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_D1 = LIOB33_X0Y5_IOB_X0Y5_I;
  assign LIOI3_SING_X0Y0_OLOGIC_X0Y0_T1 = 1'b1;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_LL2TLPRCV = 1'b0;
  assign RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y44_D = RIOB33_X43Y43_IOB_X1Y44_I;
  assign RIOI3_TBYTESRC_X43Y43_ILOGIC_X1Y43_D = RIOB33_X43Y43_IOB_X1Y43_I;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DLRSTN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPADDR8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPCLK = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPDI15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPEN = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_DRPWE = 1'b0;
  assign LIOB33_X0Y3_IOB_X0Y4_O = LIOB33_X0Y7_IOB_X0Y8_I;
  assign LIOB33_X0Y3_IOB_X0Y3_O = PCIE_BOT_X71Y115_PCIE_X0Y0_DRPRDY;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA16 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA17 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA18 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA19 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA20 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA21 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA22 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA23 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA24 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA25 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA26 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA27 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA28 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA29 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA30 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA31 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA32 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA33 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA34 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA35 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA36 = 1'b0;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_D1 = LIOB33_X0Y7_IOB_X0Y8_I;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA37 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA38 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA39 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA40 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA41 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA42 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA43 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA44 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA45 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA46 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA47 = 1'b0;
  assign LIOI3_X0Y3_OLOGIC_X0Y4_T1 = 1'b1;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA48 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA49 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA50 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA51 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA52 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA53 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA54 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA55 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA56 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA57 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA58 = 1'b0;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_D1 = PCIE_BOT_X71Y115_PCIE_X0Y0_DRPRDY;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA59 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA60 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA61 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA62 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA63 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA64 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA65 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA66 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMRXRDATA67 = 1'b0;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_D1 = RIOB33_X43Y47_IOB_X1Y47_I;
  assign LIOI3_X0Y3_OLOGIC_X0Y3_T1 = 1'b1;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y37_T1 = 1'b1;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA0 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA1 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA2 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA3 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA4 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA5 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA6 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA7 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA8 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA9 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA10 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA11 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA12 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA13 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA14 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA15 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA16 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA17 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA18 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA19 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA20 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA21 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA22 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA23 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA24 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA25 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA26 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA27 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA28 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA29 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA30 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA31 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA32 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA33 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA34 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA35 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA36 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA37 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA38 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA39 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA40 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA41 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA42 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA43 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA44 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA45 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA46 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA47 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA48 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA49 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA50 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA51 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA52 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA53 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA54 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA55 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA56 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA57 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA58 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA59 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA60 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA61 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA62 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA63 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA64 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA65 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA66 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA67 = 1'b0;
  assign PCIE_BOT_X71Y115_PCIE_X0Y0_MIMTXRDATA68 = 1'b0;
  assign RIOI3_TBYTETERM_X43Y37_OLOGIC_X1Y38_D1 = RIOB33_X43Y45_IOB_X1Y45_I;
  assign RIOB33_X43Y75_IOB_X1Y76_O = RIOB33_X43Y43_IOB_X1Y43_I;
  assign RIOB33_X43Y75_IOB_X1Y75_O = RIOB33_X43Y39_IOB_X1Y39_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_D1 = LIOB33_X0Y111_IOB_X0Y112_I;
  assign LIOI3_X0Y111_OLOGIC_X0Y111_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1 = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1 = 1'b1;
  assign LIOI3_X0Y111_ILOGIC_X0Y112_D = LIOB33_X0Y111_IOB_X0Y112_I;
  assign RIOI3_X43Y39_ILOGIC_X1Y40_D = RIOB33_X43Y39_IOB_X1Y40_I;
  assign RIOI3_X43Y39_ILOGIC_X1Y39_D = RIOB33_X43Y39_IOB_X1Y39_I;
endmodule
